`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.12.2019 07:59:36
// Design Name: 
// Module Name: simTester_verilog
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simTester_verilog();
reg CLK_100, locked, RST_IN,start_sig;
wire  completed;
localparam time t_100 = 40;

localparam integer ADDR_WIDTH = 12;
localparam integer INST_BRAM_SIZE = 2**ADDR_WIDTH;//(2**ADDR_WIDTH)
localparam integer ADDR_WIDTH_DATA_BRAM = 10;
localparam integer DATA_BRAM_SIZE = 2**ADDR_WIDTH_DATA_BRAM;//(2**ADDR_WIDTH_DATA_BRAM)
localparam integer CTRL_WIDTH = 357;
localparam integer AU_SEL_WIDTH = 5;
localparam integer BRAM_SEL_WIDTH = 5;

//This parameter = no. of BRAMS
localparam integer BRAM_LIMIT_IND_DEBUG = 8; //It indicates that BRAM contents from location 0 to BRAM_LIMIT_IND_DEBUG will be dumped for all 8 BRAMS for every cycle

//Constant array to load the A matrix
localparam integer A_size = 5892;
localparam longint A[0:5891] = '{64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc767bc81c82997, 64'hbf50f586b527553b, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbf50f586b44adc52, 64'h3fc767bc81c66fac, 64'hbd7864d9078805ad, 64'hbfc745d1745d1704, 64'h3fc767bc81c5ecca, 64'hbf50f586b408fd0b, 64'hbd7864d906ad9b68, 64'hbf50f586b32c8421, 64'h3fc767bc81c432df, 64'hbd7864d8bbbf059f, 64'hbfc745d1745d1704, 64'h3fc75e5f8dc7c993, 64'hbf488e1969eec219, 64'hbfc745d1745ddaa4, 64'hbf488e196979040c, 64'h3fc75e5f8dc7535b, 64'hbd7864d935454ad5, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4b60, 64'hbd8704e36d93dc7a, 64'hbfc745d1745d1704, 64'hbd7864d920efb5ec, 64'hbd8704e2fa09a0e9, 64'h3fc745d1745f4b60, 64'hbfc745d1745d1704, 64'hbd7864d920efb5ec, 64'h3fc745d1745f4b60, 64'hbd8704e2d324b057, 64'hbd7864d8bb51cf84, 64'hbd8704e1e81beb09, 64'h3fc745d1745f4b60, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc8169b924e1026c, 64'hbfc745d1745ddaa4, 64'hbbfe9bd2cca449db, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc75933976105d9, 64'hbf436223032b55f8, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbf436223032b55f8, 64'h3fc75933976105d9, 64'hbd7864d952e3d380, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc955503298f218e, 64'hbd7864d952e3d380, 64'hbc1304bae0f0586d, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fc745d17460474b, 64'hbd93654400792c4a, 64'hbfc745d1745ddaa4, 64'hbd32e3da3016a3ed, 64'h3fc745d1745dad9b, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc7612e1a01223a, 64'hbf4b5ca5a34823fc, 64'hbfc745d1745ddaa4, 64'hbf4b5ca5a2b82e7d, 64'h3fc7612e1a0092ad, 64'hbd7864d9376c5bc6, 64'hbfc745d1745d1704, 64'h3fc75e5f8dc447ab, 64'hbf488e19666d6e17, 64'hbd7864d8a0af0401, 64'hbfc745d1745d1704, 64'hbf488e196758ec5b, 64'h3fc75e5f8dc532b3, 64'hbd7864d8dbae6200, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbae6eadc1c86e2f2, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbae6eadb9f4153bc, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc77c75bc106647, 64'hbf5b5223d9459781, 64'hbfc745d1745ddaa4, 64'hbf5b5223d9046c5f, 64'h3fc77c75bc0fe364, 64'hbfc745d1745d1704, 64'hbd7864d9458339f9, 64'h3fc745d1745ddaa4, 64'hbca1b0c43c1a934a, 64'hbfc745d1745ddaa4, 64'hbc1fbda2dc021a17, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc75b1826022a10, 64'hbf4546b1a45032a3, 64'hbfc745d1745ddaa4, 64'hbf4546b1a407b03e, 64'h3fc75b182601e24a, 64'hbd7864d9417ef790, 64'hbfc745d1745d1704, 64'h3fc75b1826022b79, 64'hbf4546b1a450c5a3, 64'hbfc745d1745ddaa4, 64'hbf4546b1a408433d, 64'h3fc75b182601e24a, 64'hbd7864d9417ef790, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2c7cd7, 64'hbf5ad3256751484c, 64'h3fd745d5a61aff32, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca0aced851dc97a, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbc1de6740ef26f5f, 64'h3fc745d1745da3c1, 64'hbd7864d94546a2f8, 64'hbf5ad32567103494, 64'hbfc745d1745d1704, 64'h3fc77b77bf2bfb5d, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ef6ef, 64'hbd81c3c95a968962, 64'hbd74827fe4f2e1ba, 64'hbfc745d1745d1704, 64'hbd72b9312567098d, 64'h3fc745d1745e50dd, 64'hbd74827fe4f28ab0, 64'hbfc745d1745d1704, 64'h3fc745d1745f11ac, 64'hbd8566d44142127e, 64'hbd719799812dea11, 64'hbd24b4aea68a1c04, 64'h3fc745d1745da962, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61dfdecf161ab4, 64'hbc98c66deb8adaa9, 64'h3c98c66deb8adaa9, 64'h3d61dfdecf161ab4, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745dfb03, 64'hbd7468440e715093, 64'hbfc745d1745dfb03, 64'hbd7468440e715a3f, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd719777ab133f88, 64'h3ff0000000000000, 64'h3fd745d1745f26c8, 64'hbfc745d1745e15c0, 64'hbd710fb27774e48f, 64'hbfc745d1745e0a7e, 64'hbd6d120ac427d47f, 64'hbd81a0c25c277232, 64'hbd46c4a56e8c7815, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd544edbd2e8b62a, 64'h3d544edbd2e8b62a, 64'hbd65a9ce19ce2691, 64'h3d65a9ce19ce2691, 64'h3fd745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b26465de, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a935, 64'hbd719799812dea11, 64'hbd75faab2fc6ad9d, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbfc745d1745d1704, 64'hbd7864d9521f946a, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbfc745d1745d1704, 64'hbd7864d9521d5bbc, 64'h3fc745d1746079f6, 64'hbd94fd61438a8f2e, 64'hbd719799812dea11, 64'hbd3493f9ef9a9a3f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc87cf7b95f908f0, 64'hbd7864d952e2d80b, 64'hbfc745d1745d1704, 64'hbc87cf7b95f61e4a, 64'h3fc745d1745ddaa4, 64'hbd7864d952e2d80b, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8ce83533, 64'hbd7864d84b49a3cb, 64'hbc87cf797e790ba2, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'hbfc745d1745d1704, 64'hba5152ca6ad03a4b, 64'h3a5152ca6ad03a4b, 64'h3fd745d1745d1704, 64'hbddbd078fc07049d, 64'h3ddbd078fc07049d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb52298fbea1bd00, 64'h3b52298fbea1bd00, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e0c75, 64'hbf43622300319a44, 64'hbd7864d84bb6b336, 64'hbf436222fe399003, 64'h3fc75933975c149e, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1ac9, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33ad402, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b264671b, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a1a7, 64'hbd719799812dea11, 64'hbd75faab2fc6a5e0, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbfc745d1745d1704, 64'hbd7864d9521f946a, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbfc745d1745d1704, 64'hbd7864d9521d5bbc, 64'h3fc745d1746079f6, 64'hbd94fd61438a8f2e, 64'hbd719799812dea11, 64'hbd3493f9ef9a9a3f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc87cf7b95f90e02, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'hbc87cf7b95f6123f, 64'h3fc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8ce82741, 64'hbd7864d84b49a3cb, 64'hbc87cf797e790ecd, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'hbfc745d1745d1704, 64'hba51bafc9887d300, 64'h3a51bafc9887d300, 64'h3fd745d1745d1704, 64'hbddbd078fc06f886, 64'h3ddbd078fc06f886, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb52298f5674491e, 64'h3b52298f5674491e, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e0c75, 64'hbf43622300319a44, 64'hbd7864d84bb6b336, 64'hbf436222fe399003, 64'h3fc75933975c149e, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1ac9, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33ad402, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc767bc81c82997, 64'hbf50f586b527553b, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbf50f586b44adc52, 64'h3fc767bc81c66fac, 64'hbd7864d9078805ad, 64'hbfc745d1745d1704, 64'h3fc767bc81c5ecca, 64'hbf50f586b408fd0b, 64'hbd7864d906ad9b68, 64'hbf50f586b32c8421, 64'h3fc767bc81c432df, 64'hbd7864d8bbbf059f, 64'hbfc745d1745d1704, 64'h3fc75e5f8dc7c993, 64'hbf488e1969eec219, 64'hbfc745d1745ddaa4, 64'hbf488e196979040c, 64'h3fc75e5f8dc7535b, 64'hbd7864d935454ad5, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4b60, 64'hbd8704e36d944207, 64'hbfc745d1745d1704, 64'hbd7864d920f11407, 64'hbd8704e2fa0d2ff5, 64'h3fc745d1745f4b60, 64'hbfc745d1745d1704, 64'hbd7864d920f11407, 64'h3fc745d1745f4b60, 64'hbd8704e2d327744a, 64'hbd7864d8bb51cf84, 64'hbd8704e1e81b857c, 64'h3fc745d1745f4b60, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc8169b924e1026c, 64'hbfc745d1745ddaa4, 64'hbbfe9bd2cca449db, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75933976105d9, 64'hbf436223032b55f8, 64'hbd7864d952e3d380, 64'hbfc745d1745d1704, 64'hbf436223032b55f8, 64'h3fc75933976105d9, 64'hbd7864d952e3d380, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc955503298f218e, 64'hbd719799812dea11, 64'hbc1304bae0f0586d, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc22a2dc3085cbb9, 64'h3c22a2dc3085cbb9, 64'hbfc745d1745d1704, 64'hbc177b88057c8376, 64'h3c177b88057c8376, 64'h3fd745d1745d1704, 64'hbd805694f2574030, 64'h3d805694f2574030, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc8f9ac13a925d4a, 64'h3c8f9ac13a925d4a, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d17460447b, 64'hbd935230769fd6ab, 64'hbd719799812dea11, 64'hbd32d22cbe73bf2c, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc762b4c4695681, 64'hbf4ce3500b7bc7da, 64'hbd7864d938dee4ee, 64'hbf4ce3500aec6613, 64'h3fc762b4c468c6f4, 64'hbfc745d1745d1704, 64'h3fc75e5f8dc5dfcf, 64'hbf488e1968060b05, 64'hbfc745d1745ddaa4, 64'hbf488e19662f10a6, 64'h3fc75e5f8dc409bf, 64'hbd7864d8dc691fc3, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc8501bf3eb0c89d, 64'hbfc745d1745ddaa4, 64'hbc0285ef1f5121f6, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd83c04a3d1db37f, 64'h3d83c04a3d1db37f, 64'hbc7ef04364895a72, 64'h3c7ef04364895a72, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc9262d5dc729c77, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbc126511af35da74, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174ca31c7, 64'hbdeb234842dc9f4f, 64'hbd719799812dea11, 64'hbd74a7742a099eaf, 64'h3fc745d1745e49d3, 64'hbfc745d1745d1704, 64'h3fc745d17460474b, 64'hbd93654400792c4a, 64'hbfc745d1745ddaa4, 64'hbd32e3da3016a3ed, 64'h3fc745d1745dad9b, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc7612e1a01223a, 64'hbf4b5ca5a34823fc, 64'hbfc745d1745ddaa4, 64'hbf4b5ca5a2b82e7d, 64'h3fc7612e1a0092ad, 64'hbd7864d9376c5bc6, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b264671b, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a32a, 64'hbd719799812dea11, 64'hbd75faab2fc6a7cf, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbfc745d1745d1704, 64'hbd7864d9521f946a, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbfc745d1745d1704, 64'hbd7864d9521d5bbc, 64'h3fc745d1746079f6, 64'hbd94fd61438a8f2e, 64'hbd719799812dea11, 64'hbd3493f9ef9a9a3f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc87cf7b95f90e02, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'hbc87cf7b95f6123f, 64'h3fc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8ce82741, 64'hbd7864d84b49a3cb, 64'hbc87cf797e790ecd, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'hbfc745d1745d1704, 64'hba51bafc9887d300, 64'h3a51bafc9887d300, 64'h3fd745d1745d1704, 64'hbddbd078fc06fb8b, 64'h3ddbd078fc06fb8b, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb52298f5674491e, 64'h3b52298f5674491e, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e0c75, 64'hbf43622300319a44, 64'hbd7864d84bb6b336, 64'hbf436222fe399003, 64'h3fc75933975c149e, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1ac9, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33ad402, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b264671b, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a1a7, 64'hbd719799812dea11, 64'hbd75faab2fc6a5e0, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbfc745d1745d1704, 64'hbd7864d9521f946a, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbfc745d1745d1704, 64'hbd7864d9521d5bbc, 64'h3fc745d1746079f6, 64'hbd94fd61438a8f2e, 64'hbd719799812dea11, 64'hbd3493f9ef9a9a3f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc87cf7b95f90e02, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'hbc87cf7b95f6123f, 64'h3fc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8ce82741, 64'hbd7864d84b49a3cb, 64'hbc87cf797e790ecd, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'hbfc745d1745d1704, 64'hba51bafc9887d300, 64'h3a51bafc9887d300, 64'h3fd745d1745d1704, 64'hbddbd078fc06f886, 64'h3ddbd078fc06f886, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb52298f5674491e, 64'h3b52298f5674491e, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e0c75, 64'hbf43622300319a44, 64'hbd7864d84bb6b336, 64'hbf436222fe399003, 64'h3fc75933975c149e, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1ac9, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33ad402, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b264671b, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a32a, 64'hbd719799812dea11, 64'hbd75faab2fc6a7cf, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ae5ce750, 64'hbfc745d1745ddaa4, 64'hbd3cc867485320ba, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbfc745d1745d1704, 64'hbd7864d9521f946a, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbfc745d1745d1704, 64'hbd7864d9521d5bbc, 64'h3fc745d1746079f6, 64'hbd94fd61438a8f2e, 64'hbd719799812dea11, 64'hbd3493f9ef9a9a3f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee0ae3a, 64'hbd7864d91319871b, 64'hbf37e3809d9a0e98, 64'h3fc751c334aca768, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc87cf7b962d120b, 64'hbd7864d95320f7b5, 64'hbfc745d1745d1704, 64'hbc87cf7b96e28e12, 64'h3fc745d1745ddaa4, 64'hbd7864d95320f7b5, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8dd5115d, 64'hbd7864d84b49a3cb, 64'hbc87cf797ead811f, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'hbfc745d1745d1704, 64'h3ab0d9d58414687d, 64'hbab0d9d58414687d, 64'h3fd745d1745d1704, 64'hbddbd078fc06fb8b, 64'h3ddbd078fc06fb8b, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb522dd786fe7ef2, 64'h3b522dd786fe7ef2, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e0c75, 64'hbf43622300319a44, 64'hbd7864d84bb6b336, 64'hbf436222fe399003, 64'h3fc75933975c149e, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1ac9, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33ad402, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745fa40a, 64'hbd8c9bb076cf91c7, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbd1763c9b264671b, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174a320f9, 64'hbde15f254b33a32a, 64'hbd719799812dea11, 64'hbd75faab2fc6a7cf, 64'h3fc745d1745e53ad, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109ade68fa1, 64'hbfc745d1745ddaa4, 64'hbd3cc86747de0802, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc751c334ad4aa9, 64'hbf37e3809ee165f9, 64'hbfc745d1745ddaa4, 64'hbf37e3809d9ac658, 64'h3fc751c334aca768, 64'hbd7864d91319871b, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7b95f90e02, 64'hbfc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbc87cf7b95f6123f, 64'h3fc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc87cf7c8ce8269f, 64'hbd7864d952e2d23e, 64'hbc87cf797e790f6f, 64'h3fc745d1745ddaa4, 64'hbd7864d84b49a3cb, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d174617e53, 64'hbd9d21099471a475, 64'hbd719799812dea11, 64'hbd3cc8672eadb4a1, 64'h3fc745d1745db1d4, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc751c334ad5e5d, 64'hbf37e3809f08e5d1, 64'hbd7864d91319871b, 64'hbf37e3809dc2462f, 64'h3fc751c334acbb1c, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc767bc81ca60c3, 64'hbf50f586b642d03c, 64'hbd7864d9521f946a, 64'hbfc745d1745d1704, 64'hbf50f586b6409361, 64'h3fc767bc81ca5b22, 64'hbd7864d9521d5bbc, 64'hbfc745d1745d1704, 64'h3fc745d1746079f6, 64'hbd94fd6130dcb5bb, 64'hbd719799812dea11, 64'hbd3493f9dd4458e2, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hba51bafc9887d300, 64'h3a51bafc9887d300, 64'hbd15462a118bf526, 64'h3d15462a118bf526, 64'h3fd745d1745d1704, 64'hbddbd078fc06fb8b, 64'h3ddbd078fc06fb8b, 64'hbb52298f51e8387f, 64'h3b52298f51e8387f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf276434, 64'hbf5ad32564c50aa3, 64'hbd7864d9454477d5, 64'hbf5ad3256483ec1d, 64'h3fc77b77bf26e2ba, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca30c40b37740da, 64'hbd719799812dea11, 64'hbc2119fb533b629e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d174617e53, 64'hbd9d2109a6d93c7a, 64'hbfc745d1745ddaa4, 64'hbd3cc8673704ec26, 64'h3fc745d1745db1d4, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc752da1986de88, 64'hbf3a114a52090205, 64'hbfc745d1745ddaa4, 64'hbf3a114a4d3489fa, 64'h3fc752da198474b1, 64'hbd7864d87156cb39, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd92b79e9ca28724, 64'h3d92b79e9ca28724, 64'hbd85ef2b06048de3, 64'h3d85ef2b06048de3, 64'h3fd745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7593397600885, 64'hbf436223022d7375, 64'hbd7864d8cf83c829, 64'hbfc745d1745d1704, 64'hbf43622300356934, 64'h3fc75933975e0f46, 64'hbd7864d8cea9a576, 64'hbfc745d1745d1704, 64'h3fc75933975e2a03, 64'hbf436223004f4805, 64'hbd7864d84bb6b336, 64'hbf436222fe573dc4, 64'h3fc75933975c322c, 64'hbfc745d1745d1704, 64'h3fc77c75bc12a314, 64'hbf5b5223da646dcc, 64'hbfc745d1745ddaa4, 64'hbf5b5223da2340dc, 64'h3fc77c75bc122199, 64'hbd7864d9458339f9, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca1b0c38e4b1473, 64'hbfc745d1745ddaa4, 64'hbc1fbda1a33acbe5, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b793c73afb0, 64'hbf45a7c815d516dc, 64'hbd7864d930366592, 64'hbf45a7c81542384a, 64'h3fc75b793c731d52, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1746048b4, 64'hbd9375d8cd05b074, 64'hbd719799812dea11, 64'hbd3303b52f35183f, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbfc745d1745ddaa4, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbd7864d92f7b398e, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b1826021ece, 64'hbf4546b1a4446996, 64'hbd7864d92f9b5dfd, 64'hbf4546b1a3b1549c, 64'h3fc75b1826018c70, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fb7d0b12f, 64'hbd719799812dea11, 64'hbd32d22c03f5f36a, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87c9155ddd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa299f048e, 64'h3d62b1c2ff40d82e, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b6c7fe92b6, 64'h3d61e2b6c7fe92b6, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3fe1745d1746e8a0, 64'hbfc745d1745e1b62, 64'hbd704ea24540fada, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23bfb5, 64'hbd719799812dea11, 64'hbc14ce832c657224, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b688f8, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3f3f, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115ee1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcc05d, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e3053d13, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19867b1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c213a, 64'h3fc745d1745da3c1, 64'hbd7864d040a9af7b, 64'hbc6a8cff5010d1fb, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce0769, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00851, 64'hbd7864d8e3776afc, 64'hbf4484a00e1e5e26, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b68c6c43920, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd10834521ce8bf3, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce650ba2f95d2, 64'hbd719799812dea11, 64'hbd6e6d389c0e843b, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f260, 64'hbd7864d9068b4dc5, 64'hbeb46391e91120fb, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62fede, 64'hbd7864d8e315b6cb, 64'hbeb46391af34a369, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd87567afa251bdc, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106cafba9032fa, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce6788144285c, 64'hbd719799812dea11, 64'hbd6e6fbcad0e94c5, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fe3dfc9a34fe, 64'h3dd6fe3dfc9a34fe, 64'hbd5ea000a0073766, 64'h3d5ea000a0073766, 64'hbd666cac987dda0e, 64'h3d666cac987dda0e, 64'hbdd6fb887917cd77, 64'h3dd6fb887917cd77, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f80bf3a2cd316, 64'h3d7f80bf3a2cd316, 64'hbd7e007c35e53b78, 64'h3d7e007c35e53b78, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fb1bfccaf2, 64'h3d7582fb1bfccaf2, 64'hbd7e2d0a84e5774b, 64'h3d7e2d0a84e5774b, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35e94d37, 64'h3cb10b9e35e94d37, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7f01f57a92e, 64'hb529f7f01f57a92e, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df9cf, 64'hafec1bb47f3df9cf, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d6fcf0c986, 64'h3b62c2d6fcf0c986, 64'h3fd745d1745d1704, 64'hbd61dcf9ee9f136e, 64'h3d61dcf9ee9f136e, 64'hbc9a4aa0b0a6fc2c, 64'h3c9a4aa0b0a6fc2c, 64'hbc91471f29ccad6a, 64'h3c91471f29ccad6a, 64'hbe3e4b88f3083c7a, 64'h3e3e4b88f3083c7a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085790b1dcce, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564ab2, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3680b1b, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdf8d1229288, 64'hbdb7c65ac987f0e2, 64'h3db59367996233a0, 64'hbfc745d1745e5d87, 64'hbd32cd281b32fda9, 64'hbdb7d1bbd35bd060, 64'h3db59ec8a336131e, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a6471e, 64'hbfc745d1745e61c0, 64'hbd5e18a46f9d50e6, 64'hbfc745d1745e9fad, 64'h3d13ebfbce932084, 64'hbfc745d1745dea20, 64'hbd767b8bff1d827f, 64'hbfc745d1745df129, 64'hbd7598497724915c, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0a8, 64'h3c9c51d9bd23f0a8, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'hbfc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbd7864d952e46492, 64'hbd7864d84b481176, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0db040458, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fbe3233, 64'h3d4a1e6c28e04fe8, 64'h3ff0000000000000, 64'hbd92b79e90afb3af, 64'h3d92b79e90afb3af, 64'hbd6749102a1c6b53, 64'h3d6749102a1c6b53, 64'hbd8ad2076d7b5ffe, 64'h3d8ad2076d7b5ffe, 64'hbd81ac51ccec1a5a, 64'h3d81ac51ccec1a5a, 64'hbd6498d892726eda, 64'h3d6498d892726eda, 64'hbd8895908f1a877e, 64'h3d8895908f1a877e, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e97a174, 64'h3db93e221e71e432, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'h3fed1745d176b66c, 64'hbfc745d1745f18b5, 64'h3d76418c1aeefc62, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687ce6297a5, 64'h3d66e13992f3d232, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b182601fe70, 64'hbf4546b1a4243465, 64'hbfc745d1745ddaa4, 64'hbf4546b1a3911f6c, 64'h3fc75b1826016c12, 64'hbd7864d92f9b5dfd, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbd7864d92f7b398e, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fc902af8b, 64'hbd719799812dea11, 64'hbd32d22c14bb8f48, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87a94131cd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa3594c131, 64'h3d62b1c32f17ce36, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b72ec28e70, 64'h3d61e2b72ec28e70, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745e1b62, 64'hbd704ea2453ca1ad, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23c895, 64'hbd719799812dea11, 64'hbc14ce832c6577d2, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b6872b, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3ec3, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115e22, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcbf9e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e3053d13, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19867b1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c213a, 64'h3fc745d1745da3c1, 64'hbd7864d040a9af7b, 64'hbc6a8cff5010d1fb, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce019b, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00851, 64'hbd7864d8e3776afc, 64'hbf4484a00e1e5e26, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b6a0e9b7432, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108345db325a78, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58a1ec39607, 64'hbd719799812dea11, 64'hbd6e6c6aabcb6f3d, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f610, 64'hbd7864d9068b49e7, 64'hbeb46391e91117c1, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62fede, 64'hbd7864d8e315b6cb, 64'hbeb46391af34a369, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd87567afa251bdc, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106cafba9032fa, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce67881442b61, 64'hbd719799812dea11, 64'hbd6e6fbcad0e996a, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda0ba67ceba, 64'h3dd6fda0ba67ceba, 64'hbd5ea002c9e5ce91, 64'h3d5ea002c9e5ce91, 64'hbd666cac987dda0e, 64'h3d666cac987dda0e, 64'hbdd6fb887917cfe2, 64'h3dd6fb887917cfe2, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f80bf3a2cd316, 64'h3d7f80bf3a2cd316, 64'hbd7e007c35e53b78, 64'h3d7e007c35e53b78, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fca362b017, 64'h3d7582fca362b017, 64'hbd7e2d0c2a70d94e, 64'h3d7e2d0c2a70d94e, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35eb8b9f, 64'h3cb10b9e35eb8b9f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7f01f57a92e, 64'hb529f7f01f57a92e, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df8fe, 64'hafec1bb47f3df8fe, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d6fcf0c986, 64'h3b62c2d6fcf0c986, 64'h3fd745d1745d1704, 64'hbd61dcf9ff130c8c, 64'h3d61dcf9ff130c8c, 64'hbc9a4aa0b0a705ff, 64'h3c9a4aa0b0a705ff, 64'hbc91471f29ccb3c1, 64'h3c91471f29ccb3c1, 64'hbe3e4b88f309188a, 64'h3e3e4b88f309188a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085794e9ab13, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564a4f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3687ece, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdea5d4a46b4, 64'hbdb7c5bbd4239c58, 64'h3db592c8a3fddf16, 64'hbfc745d1745e5d87, 64'hbd32cd281b32fdf9, 64'hbdb7d1bbd35bd2cb, 64'h3db59ec8a3361589, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a6471e, 64'hbfc745d1745e61c0, 64'hbd5e189fa1ca92de, 64'hbfc745d1745e9fad, 64'h3d13ebfbce932084, 64'hbfc745d1745dea20, 64'hbd767b8bdc8c35e5, 64'hbfc745d1745df129, 64'hbd7598497724915c, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0f9, 64'h3c9c51d9bd23f0f9, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbd8ad207856127c9, 64'h3d8ad207856127c9, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd81ac51cd2acc0d, 64'h3d81ac51cd2acc0d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd6498d892bca433, 64'h3d6498d892bca433, 64'hbd889590a50299a2, 64'h3d889590a50299a2, 64'h3fd745d1745d1704, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d95320f9a4, 64'hbd7864d953228bf8, 64'hbd7864d84b480f87, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fc55cdd, 64'h3d4a1e6c2953024c, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e97a174, 64'h3db93e221e71e432, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176b66c, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687db45cebe, 64'h3d66e139c680b0ea, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b182601fe70, 64'hbf4546b1a4243465, 64'hbfc745d1745ddaa4, 64'hbf4546b1a3911f6c, 64'h3fc75b1826016c12, 64'hbd7864d92f9b5dfd, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbd7864d92f7b398e, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fc902af8b, 64'hbd719799812dea11, 64'hbd32d22c14bb8f48, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87a94131cd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa3594c131, 64'h3d62b1c32f17ce36, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b72ec28e70, 64'h3d61e2b72ec28e70, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745e1b62, 64'hbd704ea2453ca1ad, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23c895, 64'hbd719799812dea11, 64'hbc14ce832c6577d2, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b6872b, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3ec3, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115e22, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcbf9e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e3053d13, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19867b1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c213a, 64'h3fc745d1745da3c1, 64'hbd7864d040a9af7b, 64'hbc6a8cff5010d1fb, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce019b, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00851, 64'hbd7864d8e3776afc, 64'hbf4484a00e1e5e26, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b6a0e9b7432, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108345db325a78, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58a1ec39607, 64'hbd719799812dea11, 64'hbd6e6c6aabcb6f3d, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f610, 64'hbd7864d9068b49e7, 64'hbeb46391e91117c1, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62fede, 64'hbd7864d8e315b6cb, 64'hbeb46391af34a369, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd87567afa251bdc, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106cafba9032fa, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce67881442b61, 64'hbd719799812dea11, 64'hbd6e6fbcad0e996a, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda0ba67ceba, 64'h3dd6fda0ba67ceba, 64'hbd5ea002c9e5ce91, 64'h3d5ea002c9e5ce91, 64'hbd666cac987dda0e, 64'h3d666cac987dda0e, 64'hbdd6fb887917d030, 64'h3dd6fb887917d030, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f80bf3a2cd316, 64'h3d7f80bf3a2cd316, 64'hbd7e007c35e53b78, 64'h3d7e007c35e53b78, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fca362b017, 64'h3d7582fca362b017, 64'hbd7e2d0c2a70d94e, 64'h3d7e2d0c2a70d94e, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35eb8b9f, 64'h3cb10b9e35eb8b9f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7f01f57a92e, 64'hb529f7f01f57a92e, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df8fe, 64'hafec1bb47f3df8fe, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d6fcf0c986, 64'h3b62c2d6fcf0c986, 64'h3fd745d1745d1704, 64'hbd61dcf9ff130c8c, 64'h3d61dcf9ff130c8c, 64'hbc9a4aa0b0a705ff, 64'h3c9a4aa0b0a705ff, 64'hbc91471f29ccb3c1, 64'h3c91471f29ccb3c1, 64'hbe3e4b88f309188a, 64'h3e3e4b88f309188a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085794e9ab13, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564a4f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3687ece, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdea5d4a46b4, 64'hbdb7c5bbd4239c58, 64'h3db592c8a3fddf16, 64'hbfc745d1745e5d87, 64'hbd32cd281b32fdf9, 64'hbdb7d1bbd35bd401, 64'h3db59ec8a33616bf, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a6471e, 64'hbfc745d1745e61c0, 64'hbd5e189fa1ca92de, 64'hbfc745d1745e9fad, 64'h3d13ebfbce932084, 64'hbfc745d1745dea20, 64'hbd767b8bdc8c35e5, 64'hbfc745d1745df129, 64'hbd7598497724915c, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0f9, 64'h3c9c51d9bd23f0f9, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbd8ad207856128c1, 64'h3d8ad207856128c1, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd81ac51cd2acc0d, 64'h3d81ac51cd2acc0d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd6498d892bca433, 64'h3d6498d892bca433, 64'hbd889590a50299a2, 64'h3d889590a50299a2, 64'h3fd745d1745d1704, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbd7864d952e46492, 64'hbd7864d84b480f87, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fc55cdd, 64'h3d4a1e6c2953024c, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e979f09, 64'h3db93e221e71e1c7, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176b66c, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687db45cebe, 64'h3d66e139c680b0ea, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b182601fe70, 64'hbf4546b1a4243465, 64'hbfc745d1745ddaa4, 64'hbf4546b1a3911f6c, 64'h3fc75b1826016c12, 64'hbd7864d92f9b5dfd, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbd7864d92f7b398e, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fc902af8b, 64'hbd719799812dea11, 64'hbd32d22c14bb8f48, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87c9155ddd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa3594c131, 64'h3d62b1c32f17ce36, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b6c7fe92b6, 64'h3d61e2b6c7fe92b6, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745e1b62, 64'hbd704ea2453ca1ad, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23c895, 64'hbd719799812dea11, 64'hbc14ce832c6577d2, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b6872b, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3ec3, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115e22, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcbf9e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e3053d13, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19867b1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c213a, 64'h3fc745d1745da3c1, 64'hbd7864d040a9af7b, 64'hbc6a8cff5010d1fb, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce019b, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00851, 64'hbd7864d8e3776afc, 64'hbf4484a00e1e5e26, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b6a0e9b7432, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108345db325a78, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58a1ec39607, 64'hbd719799812dea11, 64'hbd6e6c6aabcb6f3d, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f610, 64'hbd7864d9068b49e7, 64'hbeb46391e91117c1, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62fede, 64'hbd7864d8e315b6cb, 64'hbeb46391af34a369, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd87567afa251bdc, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106cafba9032fa, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce6788144285c, 64'hbd719799812dea11, 64'hbd6e6fbcad0e958c, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda0ba67ceba, 64'h3dd6fda0ba67ceba, 64'hbd5ea002c9e5ce91, 64'h3d5ea002c9e5ce91, 64'hbd666cac987dda0e, 64'h3d666cac987dda0e, 64'hbdd6fb887917ce5f, 64'h3dd6fb887917ce5f, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f80bf3a2cd316, 64'h3d7f80bf3a2cd316, 64'hbd7e007c35e53b78, 64'h3d7e007c35e53b78, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fca362b017, 64'h3d7582fca362b017, 64'hbd7e2d0c2a70d94e, 64'h3d7e2d0c2a70d94e, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35eb74a5, 64'h3cb10b9e35eb74a5, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7f01f57a92e, 64'hb529f7f01f57a92e, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df8fe, 64'hafec1bb47f3df8fe, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d6fcf0c986, 64'h3b62c2d6fcf0c986, 64'h3fd745d1745d1704, 64'hbd61dcf9ff130c8c, 64'h3d61dcf9ff130c8c, 64'hbc9a4aa0b0a705ff, 64'h3c9a4aa0b0a705ff, 64'hbc91471f29ccb3c1, 64'h3c91471f29ccb3c1, 64'hbe3e4b88f309188a, 64'h3e3e4b88f309188a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085794e9ab13, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564a4f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3687ece, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdea5d4a46b4, 64'hbdb7c5bbd4239c58, 64'h3db592c8a3fddf16, 64'hbfc745d1745e5d87, 64'hbd32cd281b32fdf9, 64'hbdb7d1bbd35bd196, 64'h3db59ec8a3361454, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a6471e, 64'hbfc745d1745e61c0, 64'hbd5e189fa1ca92de, 64'hbfc745d1745e9fad, 64'h3d13ebfbce932084, 64'hbfc745d1745dea20, 64'hbd767b8bdc8c35e5, 64'hbfc745d1745df129, 64'hbd7598497724915c, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0f9, 64'h3c9c51d9bd23f0f9, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbd8ad207856128c1, 64'h3d8ad207856128c1, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd81ac51cd2acc0d, 64'h3d81ac51cd2acc0d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd6498d892bca433, 64'h3d6498d892bca433, 64'hbd889590a50299a2, 64'h3d889590a50299a2, 64'h3fd745d1745d1704, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbd7864d952e46492, 64'hbd7864d84b480f87, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fc55cdd, 64'h3d4a1e6c2953024c, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e97a174, 64'h3db93e221e71e432, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176b66c, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687db45cebe, 64'h3d66e139c680b0ea, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77c75bc106647, 64'hbf5b5223d9459781, 64'hbd7864d9458339f9, 64'hbf5b5223d9046c5f, 64'h3fc77c75bc0fe364, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbca1b0c43c1a934a, 64'hbd719799812dea11, 64'hbc1fbda2dc021a17, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aced851dc64f, 64'hbfc745d1745ddaa4, 64'hbc1de6740ef26cf0, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b1826022a10, 64'hbf4546b1a45032a3, 64'hbfc745d1745ddaa4, 64'hbf4546b1a407b03e, 64'h3fc75b182601e24a, 64'hbd7864d9417ef790, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc75b1826022b79, 64'hbf4546b1a450c5a3, 64'hbd7864d9417ef790, 64'hbf4546b1a408433d, 64'h3fc75b182601e24a, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c7cd7, 64'hbf5ad32567513648, 64'hbfc745d1745ddaa4, 64'hbf5ad325671017c2, 64'h3fc77b77bf2bf9f4, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ef6ef, 64'hbd81c3c95a1207e4, 64'hbfc745d1745d1704, 64'hbd74827fe4932662, 64'hbd72b93122bb1668, 64'h3fc745d1745e50dd, 64'hbfc745d1745d1704, 64'hbd74827fe492cf57, 64'h3fc745d1745f11ac, 64'hbd8566d43f5946ee, 64'hbd719799812dea11, 64'hbd24b4aea4abb4c0, 64'h3fc745d1745da962, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87a954ecca, 64'h3fd745d1745f26c8, 64'hbfc745d1745e0a7e, 64'hbd6d120ac2405c67, 64'hbd81a0c25b4bd270, 64'hbd46c4a579489f99, 64'h3ff0000000000000, 64'hbc98c66deb8ad4a3, 64'h3c98c66deb8ad4a3, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b72e5a315f, 64'h3d61e2b72e5a315f, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab133f88, 64'hbfc745d1745dfb03, 64'hbd7468440e715093, 64'h3fe1745d1746e8a0, 64'hbfc745d1745dfb03, 64'hbd7468440e715a3f, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd544edbd2e8b62a, 64'h3d544edbd2e8b62a, 64'hbd65a9ce1bec0519, 64'h3d65a9ce1bec0519, 64'h3fd745d1745d1704, 64'hbd7864d8a0af0401, 64'h3fc75e5f8dc447ab, 64'hbf488e19666d6e17, 64'hbfc745d1745d1704, 64'hbd7864d8dbae6200, 64'hbf488e196758ec5b, 64'h3fc75e5f8dc532b3, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6eadc1c86e2f2, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbae6eadb9f4153bc, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864be26827e90, 64'h3fc750009205a9e3, 64'hbf345e3b4fa0075b, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581f08a71661f, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbbf581efe3987fb5, 64'h3fc745d1745da3c1, 64'hbd7864beb4bf305f, 64'hbf345e3b522a4c40, 64'hbfc745d1745d1704, 64'h3fc750009206eefd, 64'hbfc745d1745ddaa4, 64'h3fc75a561537367e, 64'hbf4484a0d95c1418, 64'hbd7864d89cbe365f, 64'hbf4484a0d67cffe3, 64'h3fc75a56153457d7, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a562313ea04, 64'hbf4484aeb60ef3d7, 64'hbd7864d8e37803cb, 64'hbf4484aeb44d4da2, 64'h3fc75a56231227a8, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b41cf81d671, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108329844c21f4, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58943da181e, 64'hbd719799812dea11, 64'hbd6e6c69ca95b9d6, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6272fb9, 64'hbeb46392a9e19514, 64'hbd7864d89c1e7d99, 64'hbeb463913b6801da, 64'h3fc745dba62678c4, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62c5ae, 64'hbd7864d8e3164f9a, 64'hbeb46391af359e4a, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd874cbc5a13380c, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd1065d1ba21d5ee, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce64374c8d261, 64'hbd719799812dea11, 64'hbd6e6f85a6a178fa, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda00d0d829a, 64'h3dd6fda00d0d829a, 64'hbd725437cf275d49, 64'h3d725437cf275d49, 64'hbd666c8de56b95ed, 64'h3d666c8de56b95ed, 64'hbdd6fb5e7d1147a1, 64'h3dd6fb5e7d1147a1, 64'h3ff0000000000000, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae3c907f8d6c, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb641ae2960adc661, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864be264441e3, 64'h3fc745d1745ddaa4, 64'hbc6a8cd6adee374e, 64'hbfc745d1745d1704, 64'hbd7864d8e3161f3f, 64'hbc6a8d304a656b25, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c4fab83f523bae, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd7864d8a070c376, 64'h3fc745d1745ff5ab, 64'hbd90d621cd036ba5, 64'hbfc745d1745d1704, 64'hbd785e5ebd77aaad, 64'hbfc745d1745d1704, 64'hbd90cb382e4ce79d, 64'h3fc745d1745ff442, 64'hbd719799812dea11, 64'hb0c505703975e73f, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f815655a08a, 64'hbd719799812dea11, 64'hbc14ceb6f58d4861, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f46e43132d5, 64'hbd719799812dea11, 64'hbc14ce83348a78a3, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758c9cbdfe, 64'hbf5b520c1f718ad6, 64'hbd78620415fb8eb5, 64'hbfc745d1745d1704, 64'hbf5b51fe4f551c55, 64'h3fc77c7570fc84b9, 64'hbd7861f6ea364d99, 64'hbfc745d1745d1704, 64'h3fc775d719b1a46c, 64'hbf5802d2a9e5280e, 64'hbd785ec6a7938182, 64'hbf5802bdeb2bea55, 64'h3fc775d6f03431ec, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1ea4df145, 64'hbd719799812dea11, 64'hbe40ea8a629504a7, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1a48, 64'hbd719799812dea11, 64'hbe40ea8a31ff1425, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badce00cf, 64'hbf59d51cb812e810, 64'hbd7861daabaf6d6a, 64'hbfc745d1745d1704, 64'hbf59d50ef0b1a01b, 64'h3fc7797b923f3d5c, 64'hbd7861cd7ffcdfa7, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed59fd, 64'hbd785e6de9fc6aac, 64'hbf56b173ade35748, 64'h3fc773345bb9a197, 64'hbfc745d1745d1704, 64'hbe487bd31505d0e8, 64'h3e487bd31505d0e8, 64'hbeb94c1c8433da00, 64'h3eb94c1c8433da00, 64'hbeb94c1b8e514701, 64'h3eb94c1b8e514701, 64'hbe488dba9aa94264, 64'h3e488dba9aa94264, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91471eb79b9f94, 64'h3c91471eb79b9f94, 64'hbe3e68aa6ff64219, 64'h3e3e68aa6ff64219, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91474a2af10fd4, 64'h3c91474a2af10fd4, 64'hbe3e49dd98505607, 64'h3e3e49dd98505607, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f805edc1f876e, 64'h3d7f805edc1f876e, 64'hbd7df3f13bdc3d7b, 64'h3d7df3f13bdc3d7b, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hb98d208158af80c6, 64'h398d208158af80c6, 64'h3d777a5db8d7399c, 64'hbd777a5db8d7399c, 64'hb546bfa30a22edbf, 64'h3546bfa30a22edbf, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbcfc4c8f424857d3, 64'h3cfc4c8f424857d3, 64'h3fd745d1745d1704, 64'hbd61dcfa017dc633, 64'h3d61dcfa017dc633, 64'hbc9a4aa1b3be9083, 64'h3c9a4aa1b3be9083, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3d73c061f182bcc9, 64'hbd73c061f182bcc9, 64'hbaa276fc0537c216, 64'h3aa276fc0537c216, 64'h3b806f46ab30987d, 64'hbb806f46ab30987d, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'h30374a14c83b3168, 64'hb0374a14c83b3168, 64'h3fd745d1745d1704, 64'hbd88ad18100cb787, 64'h3d88ad18100cb787, 64'hbd6419c273bb8462, 64'h3d6419c273bb8462, 64'hbd89bfd288c5eec7, 64'h3d89bfd288c5eec7, 64'hbd7e2cd861b97a24, 64'h3d7e2cd861b97a24, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745e7574, 64'hbd54188ebef6ccaf, 64'hbfc745d1745eb361, 64'h3d62ea117b37dc31, 64'h3ffa2e8ba2eba536, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745e15c0, 64'hbd7108579474184e, 64'hbd6d6ae4cb477f53, 64'hbd810a1f8b5cd3f2, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30ffae9f4e7771, 64'hbdb7c5bb24f0889d, 64'h3db592c7f4cacb5b, 64'hbfc745d1745e5d87, 64'hbd333a94fcc3f5b8, 64'hbdb7d19149bc00e3, 64'h3db59e9e199643a1, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd7874328c088ac9, 64'hbd784f04d1dfe35a, 64'hbfc745d180d92512, 64'h3e38f50e05749e6b, 64'hbe410262777da977, 64'h3e4100dc71911b1e, 64'hbfc745d180b847c9, 64'h3e38b354952a1b9d, 64'hbe40d51c7b448664, 64'h3e40d396796936be, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'hbd71978e92feaf5f, 64'hbfc745d1745e19f9, 64'hbd707309eea7166b, 64'h4002e8ba2e8d1c95, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745ddaa4, 64'hbd719775a48963bc, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd5ceb546019c6cf, 64'hbd84c753e19d9f19, 64'hbfc745d1745f1cee, 64'h3d6ffc154ca40028, 64'hbfc745d1745e9fad, 64'h3d13e1f6e8514872, 64'hbfc745d1745dff3c, 64'hbd73d17734e7c309, 64'hbfc745d1745df129, 64'hbd75984d4c208c9c, 64'hbd7864be263851b9, 64'hbd7864d8e3220f69, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b38c1859, 64'hbfc745d1745ddaa4, 64'hbd719781b3c7447a, 64'hbfc745d4984e034b, 64'h3e991f7cdf6d528e, 64'hbfc745d4984de454, 64'h3e991f7be9b0f7b6, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd889591822b6454, 64'h3d889591822b6454, 64'hbd6402ad28888ec5, 64'h3d6402ad28888ec5, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd805694dd183104, 64'h3d805694dd183104, 64'hbd63c032a224bc54, 64'h3d63c032a224bc54, 64'hbc7998fde38676b9, 64'h3c7998fde38676b9, 64'hbc8b3b931fe9b2ae, 64'h3c8b3b931fe9b2ae, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbc32f54636717f2e, 64'h3c32f54636717f2e, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbde83673f4810274, 64'h3de83673f4810274, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd544edbd2ea0468, 64'h3d544edbd2ea0468, 64'hbd7b68fe378859b6, 64'h3d7b68fe378859b6, 64'h3fd745d1745d1704, 64'hbfc745d1745ddaa4, 64'hbd7197906555569b, 64'h3fed1745d176c425, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d910f5f7ac, 64'hbd7864ef255b18a5, 64'hbd719783aeb6a489, 64'hbfc745d1745e19f9, 64'hbd7079f714a85938, 64'hbfc745d1745ddaa4, 64'hbd719786b690fed2, 64'hbdb735a4c84f293f, 64'h3db502b198296bfd, 64'h3ff0000000000000, 64'hbfc745d1745e8d61, 64'hbd3f4001a8fb6602, 64'hbd876ad90718b410, 64'hbd3f3ffb43b375b0, 64'hbfc745d1745e00a4, 64'hbd738d31b1fbfecd, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176ecf6, 64'hbfc745d1745ddaa4, 64'hbd7864d8cef9d02f, 64'hbd7864d9c7b48e43, 64'hbd7864d8148e5548, 64'hbfc745d1745eb1f8, 64'h3d62b1c51226daa4, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b182601fe70, 64'hbf4546b1a4243465, 64'hbfc745d1745ddaa4, 64'hbf4546b1a3911f6c, 64'h3fc75b1826016c12, 64'hbd7864d92f9b5dfd, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbd7864d92f7b398e, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fc902af8b, 64'hbd719799812dea11, 64'hbd32d22c14bb8f48, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87c9155ddd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa3594c131, 64'h3d62b1c32f17ce36, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b6c7fe92b6, 64'h3d61e2b6c7fe92b6, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745e1b62, 64'hbd704ea2453ca1ad, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23c895, 64'hbd719799812dea11, 64'hbc14ce832c6577d2, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b6872b, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3ec3, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115e22, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcbf9e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e3053d13, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19867b1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c213a, 64'h3fc745d1745da3c1, 64'hbd7864d040a9af7b, 64'hbc6a8cff5010d1fb, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce019b, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00851, 64'hbd7864d8e3776afc, 64'hbf4484a00e1e5e26, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b6a0e9b7432, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108345db325a78, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58a1ec39607, 64'hbd719799812dea11, 64'hbd6e6c6aabcb6f3d, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f610, 64'hbd7864d9068b49e7, 64'hbeb46391e91117c1, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62fede, 64'hbd7864d8e315b6cb, 64'hbeb46391af34a369, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd87567afa251bdc, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106cafba9032fa, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce6788144285c, 64'hbd719799812dea11, 64'hbd6e6fbcad0e958c, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda0ba67cf07, 64'h3dd6fda0ba67cf07, 64'hbd5ea002c9e5ce91, 64'h3d5ea002c9e5ce91, 64'hbd666cac987dda0e, 64'h3d666cac987dda0e, 64'hbdd6fb887917ce5f, 64'h3dd6fb887917ce5f, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f80bf3a2cd316, 64'h3d7f80bf3a2cd316, 64'hbd7e007c35e53b78, 64'h3d7e007c35e53b78, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fca362b017, 64'h3d7582fca362b017, 64'hbd7e2d0c2a70d94e, 64'h3d7e2d0c2a70d94e, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35eb8b9f, 64'h3cb10b9e35eb8b9f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7f01f57a92e, 64'hb529f7f01f57a92e, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df8fe, 64'hafec1bb47f3df8fe, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d6fcf0c986, 64'h3b62c2d6fcf0c986, 64'h3fd745d1745d1704, 64'hbd61dcf9ff130c8c, 64'h3d61dcf9ff130c8c, 64'hbc9a4aa0b0a705ff, 64'h3c9a4aa0b0a705ff, 64'hbc91471f29ccb3c1, 64'h3c91471f29ccb3c1, 64'hbe3e4b88f309188a, 64'h3e3e4b88f309188a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085794e9ab13, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564a4f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3687ece, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdea5d4a46b4, 64'hbdb7c5bbd4239c58, 64'h3db592c8a3fddf16, 64'hbfc745d1745e5d87, 64'hbd32cd281b32fdf9, 64'hbdb7d1bbd35bd196, 64'h3db59ec8a3361454, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a6471e, 64'hbfc745d1745e61c0, 64'hbd5e189fa1ca92de, 64'hbfc745d1745e9fad, 64'h3d13ebfbce932084, 64'hbfc745d1745dea20, 64'hbd767b8bdc8c35e5, 64'hbfc745d1745df129, 64'hbd7598497724915c, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0f9, 64'h3c9c51d9bd23f0f9, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbd8ad207856128c1, 64'h3d8ad207856128c1, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd81ac51cd2acc0d, 64'h3d81ac51cd2acc0d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd6498d892bca433, 64'h3d6498d892bca433, 64'hbd889590a50299a2, 64'h3d889590a50299a2, 64'h3fd745d1745d1704, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d952e2d23e, 64'hbd7864d952e46492, 64'hbd7864d84b480f87, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fc55cdd, 64'h3d4a1e6c2953024c, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e97a03e, 64'h3db93e221e71e2fc, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176b66c, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687db45cebe, 64'h3d66e139c680b0ea, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d17460474b, 64'hbd9365446d0a8a40, 64'hbd719799812dea11, 64'hbd32e3da99f6b122, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7612e1a0024e7, 64'hbf4b5ca5a249ef55, 64'hbd7864d9376c5bc6, 64'hbf4b5ca5a1b9f9d6, 64'h3fc7612e19ff93f1, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbca0aceda0c3c567, 64'hbfc745d1745ddaa4, 64'hbc1de67440b02c1c, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc75b182601fe70, 64'hbf4546b1a4243465, 64'hbfc745d1745ddaa4, 64'hbf4546b1a3911f6c, 64'h3fc75b1826016c12, 64'hbd7864d92f9b5dfd, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8b774ead95fc25, 64'hbd7864d92f7b398e, 64'hbc8b774e3477fb4d, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'h3fc77b77bf2c1d24, 64'hbf5ad3256721a659, 64'hbfc745d1745ddaa4, 64'hbf5ad32566e087d3, 64'h3fc77b77bf2b9ba9, 64'hbd7864d9454477d5, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc77b77bf2d1eb0, 64'hbf5ad32567a1f066, 64'hbfc745d1745d1704, 64'hbd7864d95271bbda, 64'hbf5ad325679fce90, 64'h3fc77b77bf2d1a78, 64'hbfc745d1745d1704, 64'hbd7864d9526fb199, 64'h3fc745d17460447b, 64'hbd93522fc902af8b, 64'hbd719799812dea11, 64'hbd32d22c14bb8f48, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745e15c0, 64'hbd710e87c9155ddd, 64'h3fd745d1745f45bf, 64'hbfc745d1745ddc0d, 64'hbd7827652495d3d6, 64'hbd89aaaa3594c131, 64'h3d62b1c32f17ce36, 64'h3ff0000000000000, 64'hbc98c66e14be4f0c, 64'h3c98c66e14be4f0c, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b6c7fe92b6, 64'h3d61e2b6c7fe92b6, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745ddaa4, 64'hbd719777ab130805, 64'hbfc745d1745e1b62, 64'hbd704ea2453ca1ad, 64'h3fe1745d1746e8a0, 64'hbfc745d1745ddaa4, 64'hbd7864d92f7afba8, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbb2683a044d6ff7d, 64'h3b2683a044d6ff7d, 64'hbd12b9b8d8cf6abe, 64'h3d12b9b8d8cf6abe, 64'h3fd745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581d274e53b0e, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbbf581d1ce0d3c06, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e25bb375, 64'h3fc7500092407ccc, 64'hbf345e3bc544f073, 64'hbfc745d1745d1704, 64'hbd7864d8709a82de, 64'hbf345e3bc7cf34a0, 64'h3fc750009241c1e6, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbae6f7f3f4d4bbea, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd785ea5b4064c81, 64'h3fc75e5f74fa7cb1, 64'hbf488e009ca204ca, 64'hbfc745d1745d1704, 64'hbd785ea5eecef080, 64'hbfc745d1745d1704, 64'hbf488e009d8d8255, 64'h3fc75e5f74fb67ba, 64'hbd719799812dea11, 64'hbae6f7f377497772, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f477e23c895, 64'hbd719799812dea11, 64'hbc14ce832c6577d2, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f490d358dd5, 64'hbd719799812dea11, 64'hbc14ce8523a8b9a0, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758d2b0643, 64'hbf5b520c6695f8f9, 64'hbd786203edf23d30, 64'hbfc745d1745d1704, 64'hbf5b51fe95b6872b, 64'h3fc77c7571894726, 64'hbd7861f6c172dcee, 64'hbfc745d1745d1704, 64'h3fc775d719ac95a3, 64'hbf5802d2a75d82bd, 64'hbd785ec651cc2968, 64'hbf5802bde77ea0bb, 64'h3fc775d6f02cd6db, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1e923490c, 64'hbd719799812dea11, 64'hbe40ea8a6265dc65, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1870, 64'hbd719799812dea11, 64'hbe40ea8a31ff13ac, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badc8dce9, 64'hbf59d51cb5817abe, 64'hbd7861daabaee036, 64'hbfc745d1745d1704, 64'hbf59d50eee202b94, 64'h3fc7797b923a1adf, 64'hbd7861cd7ffc5084, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed5495, 64'hbd785e6de9fb9209, 64'hbf56b173ade34e46, 64'h3fc773345bb9a02f, 64'hbfc745d1745d1704, 64'hbe487d2da519982f, 64'h3e487d2da519982f, 64'hbeb94c1c8345308a, 64'h3eb94c1c8345308a, 64'hbeb94c1b8e514529, 64'h3eb94c1b8e514529, 64'hbe488dba9cc3e521, 64'h3e488dba9cc3e521, 64'h3ff0000000000000, 64'hbd785ea5b3c847ed, 64'h3fc745d1745ff442, 64'hbd90cde2477eacac, 64'hbfc745d1745d1704, 64'hbd785e6757716ee8, 64'hbd90cd791cec3ec3, 64'h3fc745d1745ff442, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c504a78c115e22, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb0c5050f09fcbf9e, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864d7e21d74d9, 64'h3fc745d1745ddaa4, 64'hbc6a8d18e302d276, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae37c19a0cb5, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hb641ae3d3b5c1ed1, 64'h3fc745d1745da3c1, 64'hbd7864d040abfb80, 64'hbc6a8cff50161e5e, 64'hbfc745d1745d1704, 64'h3fc745d1745ddaa4, 64'hbfc745d1745ddaa4, 64'h3fc75a5614fc1a65, 64'hbf4484a09e409d40, 64'hbd7864d906ce019b, 64'hbf4484a09d0d8fc8, 64'h3fc75a5614fae797, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a56146dba34, 64'hbf4484a00fe00db9, 64'hbd7864d8e379b702, 64'hbf4484a00e1e6cec, 64'h3fc75a56146bf940, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b6a0e9b7432, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108345db325a78, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58a1ec39607, 64'hbd719799812dea11, 64'hbd6e6c6aabcb6f3d, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6271c05, 64'hbeb463928225f610, 64'hbd7864d9068b49e7, 64'hbeb46391e91117c1, 64'h3fc745dba626ce9d, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f622359, 64'hbd7864d8e31802d1, 64'hbeb46391af38647d, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd8755ee8e94e595, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd106c608c9338c2, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174981c98, 64'hbddd3c9539b550b3, 64'hbd719799812dea11, 64'hbd6ec90cbc0c408e, 64'h3fc745d1745e1f9a, 64'hbfc745d1745d1704, 64'hbdd6fda0ba67ceba, 64'h3dd6fda0ba67ceba, 64'hbd5ea002c9e5ce91, 64'h3d5ea002c9e5ce91, 64'hbd666c367c1a04a4, 64'h3d666c367c1a04a4, 64'hbdd73faee179f173, 64'h3dd73faee179f173, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f8019566b1bad, 64'h3d7f8019566b1bad, 64'hbd7dffc794bb79c7, 64'h3d7dffc794bb79c7, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7582fca362b017, 64'h3d7582fca362b017, 64'hbd7e2d0c2a70d94e, 64'h3d7e2d0c2a70d94e, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91472052bf7e76, 64'h3c91472052bf7e76, 64'hbe3e68aa7f9738eb, 64'h3e3e68aa7f9738eb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d777a5dc1bdfd61, 64'hbd777a5dc1bdfd61, 64'hb98d30b03e6ce3da, 64'h398d30b03e6ce3da, 64'hbcb10b9e35ebf29e, 64'h3cb10b9e35ebf29e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3529f7e84b4e246f, 64'hb529f7e84b4e246f, 64'h3fd745d1745d1704, 64'hbd88ad189a58d6b3, 64'h3d88ad189a58d6b3, 64'hbd6419c25a300408, 64'h3d6419c25a300408, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276e28596c4af, 64'h3aa276e28596c4af, 64'h3d73c03de4303a10, 64'hbd73c03de4303a10, 64'h2fec1bb47f3df8fe, 64'hafec1bb47f3df8fe, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'hbb62c2d1551f0731, 64'h3b62c2d1551f0731, 64'h3fd745d1745d1704, 64'hbd61dcf9ff130c8c, 64'h3d61dcf9ff130c8c, 64'hbc9a4aa0b0a705ff, 64'h3c9a4aa0b0a705ff, 64'hbc91471f29ccb3c1, 64'h3c91471f29ccb3c1, 64'hbe3e4b88f309188a, 64'h3e3e4b88f309188a, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'hbfc745d1745f18b5, 64'h3d76418c343c9d4b, 64'hbfc745d1745e15c0, 64'hbd71085794e9ab13, 64'h3ffa2e8ba2eb9e2c, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbfc745d1745eb361, 64'h3d62ea12a9564a4f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbd6d5e6af1914502, 64'hbd81070b15064d40, 64'hbfc745d180d9d4fe, 64'h3e38f66eb3687ece, 64'hbe4103532e37bde5, 64'h3e4101cd284f2406, 64'hbfc745d180b847c9, 64'h3e38b3549d7272d6, 64'hbe40d51c7cb59b43, 64'h3e40d3967ada4b61, 64'hbd785f39a42e9f80, 64'hbd785dd3670b1754, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30fdea5d4a46b4, 64'hbdb7c5bbd4239c58, 64'h3db592c8a3fddf16, 64'hbfc745d1745e5d87, 64'hbd32d357af1e50c3, 64'hbdb816ca931ff4c2, 64'h3db5e3d762fa3780, 64'h3ff0000000000000, 64'hbfc745d1745ee60b, 64'h3d6208ac7e646897, 64'hbfc745d1745ddaa4, 64'hbd719775a48ac0df, 64'h4002e8ba2e8d1f38, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbfc745d1745e19f9, 64'hbd707309f1c80bd7, 64'hbd5cebb82929e3a8, 64'hbd84c7612455ddbd, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b3c6a57b, 64'hbfc745d1745ddaa4, 64'hbd719781b3c514b2, 64'hbfc745d4984e034b, 64'h3e991f7cde7ecf18, 64'hbfc745d4984de454, 64'h3e991f7be9b0f580, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd7864d7e220dd35, 64'hbd7864d040a89324, 64'hbfc745d1745e61c0, 64'hbd5e189fa1ca92de, 64'hbfc745d1745e9fad, 64'h3d13cb74c2f9ed02, 64'hbfc745d1745dea20, 64'hbd767b8bdc8c35e5, 64'hbfc745d1745df129, 64'hbd759858354e9671, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd61e2b733f11cba, 64'h3d61e2b733f11cba, 64'hbc9c51d9bd23f0f9, 64'h3c9c51d9bd23f0f9, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbd8272016ef55f28, 64'h3d8272016ef55f28, 64'hbd92b79ea1107ac3, 64'h3d92b79ea1107ac3, 64'hbd6749102a62ef33, 64'h3d6749102a62ef33, 64'hbd81ac51ca8c0ff7, 64'h3d81ac51ca8c0ff7, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbd8ad207856127c9, 64'h3d8ad207856127c9, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd81ac51cd2acc0d, 64'h3d81ac51cd2acc0d, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd6498d892bca433, 64'h3d6498d892bca433, 64'hbd889590a50299a2, 64'h3d889590a50299a2, 64'h3fd745d1745d1704, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafdb78a, 64'h3fed1745d176faae, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd7864d952e2d80b, 64'hbd7864d952e46a60, 64'hbd7864d84b480f87, 64'hbfc745d1745ddaa4, 64'hbd719772ef5f1d6d, 64'hbfc745d1745eb79a, 64'h3d4a1e682681eeb6, 64'hbd8a06bf4fc55cdd, 64'h3d4a1e6c2953024c, 64'h3ff0000000000000, 64'hbfc745d1745e79ad, 64'h3d42f1ab3de7541d, 64'hbdbb71154e97ab20, 64'h3db93e221e71edde, 64'hbfc745d1745f18b5, 64'h3d76418c3dac8a12, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176b66c, 64'hbfc745d1745ddc0d, 64'hbd782a6884122275, 64'hbd8ab687db45cebe, 64'h3d66e139c680b0ea, 64'hbfc745d1745e15c0, 64'hbd710e87a84665c8, 64'h3ff0000000000000, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'hbd648fd74e1a81b7, 64'h3d648fd74e1a81b7, 64'hbd88cf672e8cdec3, 64'h3d88cf672e8cdec3, 64'h3ff0000000000000, 64'hbd7864be26827e90, 64'h3fc750009205a9e3, 64'hbf345e3b4fa0075b, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hbbf581f08a71661f, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbbf581efe3987fb5, 64'h3fc745d1745da3c1, 64'hbd7864beb4bf305f, 64'hbf345e3b522a4c40, 64'hbfc745d1745d1704, 64'h3fc750009206eefd, 64'hbfc745d1745ddaa4, 64'h3fc75a561537367e, 64'hbf4484a0d95c1418, 64'hbd7864d89cbe365f, 64'hbf4484a0d67cffe3, 64'h3fc75a56153457d7, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75a562313ea04, 64'hbf4484aeb60ef3d7, 64'hbd7864d8e37803cb, 64'hbf4484aeb44d4da2, 64'h3fc75a56231227a8, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f5269, 64'hbd877b41cf81d671, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd108329844c21f4, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174976f7d, 64'hbddce58943da181e, 64'hbd719799812dea11, 64'hbd6e6c69ca95b9d6, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745dba6272fb9, 64'hbeb46392a9e19514, 64'hbd7864d89c1e7d99, 64'hbeb463913b6801da, 64'h3fc745dba62678c4, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745dba62721a6, 64'hbeb463928f62c5ae, 64'hbd7864d8e3164f9a, 64'hbeb46391af359e4a, 64'h3fc745dba626b278, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745f4f99, 64'hbd874cbc5a13380c, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbd1065d1ba21d5ee, 64'h3fc745d1745da692, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d1749770e5, 64'hbddce64374c8cf5c, 64'hbd719799812dea11, 64'hbd6e6f85a6a173f3, 64'h3fc745d1745e1e32, 64'hbfc745d1745d1704, 64'hbdd6fda00d0d829a, 64'h3dd6fda00d0d829a, 64'hbd725437cf275d49, 64'h3d725437cf275d49, 64'hbd666c8de56b95ed, 64'h3d666c8de56b95ed, 64'hbdd6fb5e7d11449b, 64'h3dd6fb5e7d11449b, 64'h3ff0000000000000, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb641ae3c907f8d6c, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'hb641ae2960adc661, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd7864be264441e3, 64'h3fc745d1745ddaa4, 64'hbc6a8cd6adee374e, 64'hbfc745d1745d1704, 64'hbd7864d8e3161f3f, 64'hbc6a8d304a656b25, 64'h3fc745d1745ddaa4, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc76f9565ad1a48, 64'hbf54e1f8a79fa890, 64'hbd7864d9416d01c6, 64'hbf54e1f8a75f80d6, 64'h3fc76f9565ac98ce, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc994cca0591407e, 64'hbd719799812dea11, 64'hbc169b72502957f1, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbd719799812dea11, 64'h3fc745d1745da3c1, 64'hb0c4fab83f523bae, 64'hbfc745d1745d1704, 64'h3fd745fb65c828cb, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbee4f8b588e368f1, 64'hbd7864d8a070c376, 64'h3fc745d1745ff5ab, 64'hbd90d621cd036ba5, 64'hbfc745d1745d1704, 64'hbd785e5ebd77aaad, 64'hbfc745d1745d1704, 64'hbd90cb382e4ce79d, 64'h3fc745d1745ff442, 64'hbd719799812dea11, 64'hb0c505703975e73f, 64'hbfc745d1745d1704, 64'h3fc745d1745da3c1, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f815655a08a, 64'hbd719799812dea11, 64'hbc14ceb6f58d4861, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc974f46e43132d5, 64'hbd719799812dea11, 64'hbc14ce83348a78a3, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc77c758c9cbdfe, 64'hbf5b520c1f718ad6, 64'hbd78620415fb8eb5, 64'hbfc745d1745d1704, 64'hbf5b51fe4f551c55, 64'h3fc77c7570fc84b9, 64'hbd7861f6ea364d99, 64'hbfc745d1745d1704, 64'h3fc775d719b1a46c, 64'hbf5802d2a9e5280e, 64'hbd785ec6a7938182, 64'hbf5802bdeb2bea55, 64'h3fc775d6f03431ec, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745e14f46cf9b, 64'hbebfb5d1ea4df145, 64'hbd719799812dea11, 64'hbe40ea8a629504a7, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'h3fc745e14f463633, 64'hbebfb5d0b69b1a48, 64'hbd719799812dea11, 64'hbe40ea8a31ff1425, 64'h3fc745d185482e81, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc7797badce00cf, 64'hbf59d51cb812e810, 64'hbd7861daabaf6d6a, 64'hbfc745d1745d1704, 64'hbf59d50ef0b1a01b, 64'h3fc7797b923f3d5c, 64'hbd7861cd7ffcdfa7, 64'hbfc745d1745d1704, 64'h3fc77334851bb4c5, 64'hbf56b1885eed59fd, 64'hbd785e6de9fc6aac, 64'hbf56b173ade35748, 64'h3fc773345bb9a197, 64'hbfc745d1745d1704, 64'hbe487bd31505d0e8, 64'h3e487bd31505d0e8, 64'hbeb94c1c8433da00, 64'h3eb94c1c8433da00, 64'hbeb94c1b8e514701, 64'h3eb94c1b8e514701, 64'hbe488dba9aa94264, 64'h3e488dba9aa94264, 64'h3ff0000000000000, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91471eb79b9f94, 64'h3c91471eb79b9f94, 64'hbe3e68aa6ff64219, 64'h3e3e68aa6ff64219, 64'h3fed1745d1745d1f, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc91474a2af10fd4, 64'h3c91474a2af10fd4, 64'hbe3e49dd98505607, 64'h3e3e49dd98505607, 64'h3fe745d1745d175e, 64'hbd61dcfa017dc633, 64'h3d61dcfa017dc633, 64'hbc9a4aa1b3be9083, 64'h3c9a4aa1b3be9083, 64'hbee4f8b588e368f1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe174720ffb5a81, 64'hb98d208158af80c6, 64'h398d208158af80c6, 64'h3d777a5db8d7399c, 64'hbd777a5db8d7399c, 64'hb546bfa30a22edbf, 64'h3546bfa30a22edbf, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbcfc4c8f42485a4c, 64'h3cfc4c8f42485a4c, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd7f805edc1f876e, 64'h3d7f805edc1f876e, 64'hbd7df3f13bdc3d7b, 64'h3d7df3f13bdc3d7b, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'h3d73c061f182bcc9, 64'hbd73c061f182bcc9, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbaa276fc0537c216, 64'h3aa276fc0537c216, 64'h3b806f46ab30987d, 64'hbb806f46ab30987d, 64'hbd623c645875fc25, 64'h3d623c645875fc25, 64'hbc92c363a24925eb, 64'h3c92c363a24925eb, 64'h30374a14c83b3168, 64'hb0374a14c83b3168, 64'h3fd745d1745d1704, 64'hbd88ad18100cb787, 64'h3d88ad18100cb787, 64'hbd6419c273bb8462, 64'h3d6419c273bb8462, 64'hbd89bfd288c5eec7, 64'h3d89bfd288c5eec7, 64'hbd7e2cd861b97a24, 64'h3d7e2cd861b97a24, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe1745d1745d19d, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc9262d5dc72b255, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'hbc126511af35ddb3, 64'h3fc745d1745da3c1, 64'hbd719799812dea11, 64'hbfc745d1745d1704, 64'h3fc745d174ca31c7, 64'hbdeb234842c2e42c, 64'hbd719799812dea11, 64'hbd74a77429f627f9, 64'h3fc745d1745e49d3, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d17460447b, 64'hbd935230769fd6ab, 64'hbd719799812dea11, 64'hbd32d22cbe73bf2c, 64'h3fc745d1745dad9b, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc762b4c4695681, 64'hbf4ce3500b7bc7da, 64'hbd7864d938dee4ee, 64'hbf4ce3500aec6613, 64'h3fc762b4c468c6f4, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc75e5f8dc5dfcf, 64'hbf488e1968060b05, 64'hbd7864d8dc691fc3, 64'hbf488e19662f10a6, 64'h3fc75e5f8dc409bf, 64'hbfc745d1745d1704, 64'hbfc745d1745ddaa4, 64'h3fc745d1745ddaa4, 64'hbc8501bf3eb0c89d, 64'hbd719799812dea11, 64'hbc0285ef1f5121f6, 64'h3fc745d1745da3c1, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd83c04a3d1db37f, 64'h3d83c04a3d1db37f, 64'hbc7ef04364895a72, 64'h3c7ef04364895a72, 64'h3fd745d1745d1704, 64'hbfc745d1745eb361, 64'h3d62ea117b37dc31, 64'hbd6d6ae4cb477f53, 64'hbd810a1f8b5cd3f2, 64'hbfc745d1745e15c0, 64'hbd7108579474184e, 64'h3ffa2e8ba2eba536, 64'hbfc745d1745eb361, 64'h3d62e18005b79168, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e5eef, 64'hbd30ffae9f4e7771, 64'hbdb7c5bb24f0889d, 64'h3db592c7f4cacb5b, 64'hbfc745d1745e5d87, 64'hbd333a94fcc3f568, 64'hbdb7d19149bbfd43, 64'h3db59e9e19964001, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745e1188, 64'hbd717955b8e16ec5, 64'hbd7874328c088ac9, 64'hbd784f04d1dfe35a, 64'hbfc745d180d92512, 64'h3e38f50e05749e6b, 64'hbe410262777da977, 64'h3e4100dc71911b1e, 64'hbfc745d180b847c9, 64'h3e38b354952a1b9d, 64'hbe40d51c7b448664, 64'h3e40d396796936be, 64'hbfc745d1745e7574, 64'hbd54188ebef6ccaf, 64'h3ff0000000000000, 64'hbfc745d1745e19f9, 64'hbd707309eea7166b, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719775a48963bc, 64'h4002e8ba2e8d1c95, 64'hbfc745d1745e1b62, 64'hbd7050f5245b9c89, 64'hbd5ceb546019c6cf, 64'hbd84c753e19d9f19, 64'hbfc745d1745f1cee, 64'h3d6ffc154ca40028, 64'hbfc745d1745e9fad, 64'h3d13e1f6e8514872, 64'hbfc745d1745dff3c, 64'hbd73d17734e7c309, 64'hbfc745d1745df129, 64'hbd75984d4c208c9c, 64'hbd7864be263851b9, 64'hbd7864d8e3220f69, 64'hbfc745d1745ddaa4, 64'hbd71977fb602262f, 64'hbd719799812dea11, 64'hbd719799812dea11, 64'hbfc745d1745ddaa4, 64'hbd719781b38c1859, 64'hbfc745d1745ddaa4, 64'hbd719781b3c7447a, 64'hbfc745d4984e034b, 64'h3e991f7cdf6d528e, 64'hbfc745d4984de454, 64'h3e991f7be9b0f7b6, 64'hbfc745d1745ddaa4, 64'hbd71978e92feaf5f, 64'h3ff0000000000000, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'h3fe745d1745d175e, 64'hbfc745d1745d1704, 64'hbc22a35ed0bca9ce, 64'h3c22a35ed0bca9ce, 64'hbfc745d1745d1704, 64'hbc177b88057c8376, 64'h3c177b88057c8376, 64'h3fd745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbd889591822b6454, 64'h3d889591822b6454, 64'hbd6402ad28888ec5, 64'h3d6402ad28888ec5, 64'h3fe745d1745d175e, 64'hbd805694f2574030, 64'h3d805694f2574030, 64'hbfc745d1745d1704, 64'hbc8f9ac13a925d4a, 64'h3c8f9ac13a925d4a, 64'hbfc745d1745d1704, 64'h3fd745d1745d1704, 64'hbd805694dd183104, 64'h3d805694dd183104, 64'hbd63c032a224bc54, 64'h3d63c032a224bc54, 64'hbc7998fde38676b9, 64'h3c7998fde38676b9, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbc8b3b931fe9d301, 64'h3c8b3b931fe9d301, 64'h3fd745d1745d1704, 64'hbd92b79ea15c9e08, 64'h3d92b79ea15c9e08, 64'hbc32f504e6560e84, 64'h3c32f504e6560e84, 64'hbd6749102a643740, 64'h3d6749102a643740, 64'hbd544edbd2ea0468, 64'h3d544edbd2ea0468, 64'hbd7b68fe39f378b8, 64'h3d7b68fe39f378b8, 64'hbfc745d1745d1704, 64'hbfc745d1745d1704, 64'hbde83673f46a16a1, 64'h3de83673f46a16a1, 64'h3fd745d1745d1704, 64'hbfc745d1745e8d61, 64'hbd3f4001a8fb6602, 64'hbd876ad90718b410, 64'hbd3f3ffb43b375b0, 64'hbfc745d1745e00a4, 64'hbd738d31b1fbfecd, 64'hbfc745d1745f18b5, 64'h3d76418c3e4e0966, 64'h3fed1745d176ecf6, 64'hbfc745d1745ddaa4, 64'hbd7864d8cef63399, 64'hbd7864d9c7b0f1ad, 64'hbd7864d8149093c3, 64'hbfc745d1745eb1f8, 64'h3d62b1c51226daa4, 64'h3ff0000000000000, 64'hbfc745d1745ddaa4, 64'hbd7197906555569b, 64'hbfc745d1745ddaa4, 64'hbd7864d910f5f7ac, 64'hbd7864ef255b18a5, 64'hbd719783aeb6a489, 64'h3fed1745d176c425, 64'hbfc745d1745e2103, 64'hbd6f3ec0dafd9a23, 64'hbfc745d1745ddaa4, 64'hbd719786b690fed2, 64'hbdb735a4c839ea4a, 64'h3db502b198142d07, 64'hbfc745d1745e19f9, 64'hbd7079f714a85938, 64'h3ff0000000000000};
localparam integer A_BRAMInd[0:5891] = '{0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 0, 1, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 4, 5, 0, 2, 3, 6, 0, 1, 2, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 5, 6, 1, 3, 4, 7, 1, 2, 3, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 6, 7, 2, 4, 5, 0, 2, 3, 4, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 7, 0, 3, 5, 6, 1, 3, 4, 5, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 0, 1, 4, 6, 7, 2, 4, 5, 6, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 1, 2, 5, 7, 0, 3, 5, 6, 7, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 0, 1, 4, 6, 7, 0, 1, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 7, 1, 2, 3, 4, 6, 7, 3, 5, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 4, 6, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 6, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 3, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 2, 3, 6, 0, 2, 3, 4, 5, 1, 5, 7, 1, 2, 3, 4, 7, 0, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 1, 5, 6, 7, 0, 2, 5, 6, 7, 2, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 3, 7, 0, 1, 2, 5, 6, 7, 0, 3, 4, 5, 7, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 5, 6, 1, 2, 6, 1, 2, 5, 6, 7, 0, 4, 5, 0, 1, 4, 6, 7, 2, 3, 4, 5, 6, 0, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 3, 5, 6, 7, 0, 6, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 7, 1, 2, 3, 4, 5, 6, 2, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 3, 4, 5, 7, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 6, 1, 2, 5, 7, 1, 2, 3, 4, 0, 4, 6, 0, 1, 2, 3, 6, 7, 5, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 0, 4, 5, 6, 7, 1, 4, 5, 6, 1, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 2, 6, 7, 0, 1, 4, 5, 6, 7, 2, 3, 4, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 0, 1, 5, 0, 2, 3, 4, 5, 6, 7, 1, 5, 0, 1, 4, 5, 7, 0, 3, 4, 7, 0, 4, 6, 7, 1, 2, 3, 4, 6, 7, 0, 2, 4, 5, 7, 0, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 4, 5, 6, 7, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 3, 4, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 5, 7, 0, 1, 2, 3, 4, 0, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 0, 1, 3, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 7, 0, 3, 5, 7, 0, 1, 2, 6, 2, 4, 6, 7, 0, 1, 4, 5, 3, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 6, 2, 3, 4, 5, 7, 2, 3, 4, 7, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 0, 4, 5, 6, 7, 2, 3, 4, 5, 0, 1, 2, 4, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 6, 7, 3, 6, 0, 1, 2, 3, 4, 5, 7, 3, 6, 7, 2, 3, 5, 6, 1, 2, 5, 6, 2, 4, 5, 7, 0, 1, 2, 4, 5, 6, 0, 2, 3, 5, 6, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 7, 0, 2, 3, 4, 5, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 2, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 3, 5, 6, 7, 0, 1, 2, 6, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 5, 6, 7, 1, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 0, 1, 3, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 5, 6, 1, 3, 5, 6, 7, 0, 4, 0, 2, 4, 5, 6, 7, 2, 3, 1, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 4, 0, 1, 2, 3, 5, 0, 1, 2, 5, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 6, 2, 3, 4, 5, 0, 1, 2, 3, 6, 7, 0, 2, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 0, 1, 4, 5, 1, 4, 6, 7, 0, 1, 2, 3, 5, 1, 4, 5, 0, 1, 3, 4, 7, 0, 3, 4, 0, 2, 3, 5, 6, 7, 0, 2, 3, 4, 6, 0, 1, 3, 4, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 5, 6, 0, 1, 2, 3, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 3, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 0, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 1, 3, 4, 5, 6, 7, 0, 4, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 3, 4, 5, 7, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 5, 6, 7, 1, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 0, 3, 4, 7, 1, 3, 4, 5, 6, 2, 6, 0, 2, 3, 4, 5, 0, 1, 7, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 2, 6, 7, 0, 1, 3, 6, 7, 0, 3, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 4, 0, 1, 2, 3, 6, 7, 0, 1, 4, 5, 6, 0, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 6, 7, 2, 3, 7, 2, 4, 5, 6, 7, 0, 1, 3, 7, 2, 3, 6, 7, 1, 2, 5, 6, 1, 2, 6, 0, 1, 3, 4, 5, 6, 0, 1, 2, 4, 6, 7, 1, 2, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 3, 4, 6, 7, 0, 1, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 7, 1, 2, 3, 4, 5, 6, 2, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 3, 4, 5, 7, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 6, 1, 2, 5, 7, 1, 2, 3, 4, 0, 4, 6, 0, 1, 2, 3, 6, 7, 5, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 0, 4, 5, 6, 7, 1, 4, 5, 6, 1, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 2, 6, 7, 0, 1, 4, 5, 6, 7, 2, 3, 4, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 5, 0, 1, 5, 0, 2, 3, 4, 5, 6, 7, 1, 5, 0, 1, 4, 5, 7, 0, 3, 4, 7, 0, 4, 6, 7, 1, 2, 3, 4, 6, 7, 0, 2, 4, 5, 7, 0, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 4, 5, 6, 7, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 2, 3, 4, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 5, 7, 0, 1, 2, 3, 4, 0, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 0, 1, 3, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 7, 0, 3, 5, 7, 0, 1, 2, 6, 2, 4, 6, 7, 0, 1, 4, 5, 3, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 6, 2, 3, 4, 5, 7, 2, 3, 4, 7, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 0, 4, 5, 6, 7, 2, 3, 4, 5, 0, 1, 2, 4, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 2, 3, 6, 7, 3, 6, 0, 1, 2, 3, 4, 5, 7, 3, 6, 7, 2, 3, 5, 6, 1, 2, 5, 6, 2, 4, 5, 7, 0, 1, 2, 4, 5, 6, 0, 2, 3, 5, 6, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 7, 0, 2, 3, 4, 5, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 7, 0, 1, 3, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 6, 7, 0, 1, 2, 3, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 1, 2, 3, 5, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 0, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 4, 7, 0, 3, 5, 7, 0, 1, 2, 6, 2, 3, 4, 5, 1, 4, 5, 6, 0, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 3, 7, 1, 5, 6, 7, 0, 3, 4, 3, 6, 7, 0, 2, 3, 4, 6, 7, 0, 1, 2, 3, 4, 5, 4, 7, 0, 1, 2, 5, 6, 7, 0, 3, 4, 5, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 5, 6, 7, 0, 1, 2, 4, 5, 6, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 5, 6, 3, 4, 5, 7, 1, 2, 5, 6, 7, 3, 5, 7, 0, 2, 3, 4, 5, 6, 1, 3, 4, 5, 7, 0, 2, 4, 6, 7, 2, 3, 5, 6, 0, 1, 4, 5, 2, 3, 4, 6, 7, 0, 1, 2, 3, 5, 6, 0, 2, 4, 5, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 5};
localparam integer A_BRAMAddr[0:5891] = '{0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 48, 48, 48, 48, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 52, 52, 52, 52, 53, 53, 53, 53, 53, 53, 53, 53, 54, 54, 54, 54, 54, 54, 54, 54, 55, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 56, 56, 56, 56, 57, 57, 57, 57, 57, 57, 58, 58, 58, 58, 58, 58, 58, 58, 59, 59, 59, 59, 59, 59, 59, 59, 60, 60, 60, 60, 60, 60, 60, 60, 61, 61, 61, 61, 61, 61, 61, 62, 62, 62, 62, 62, 62, 62, 63, 63, 63, 63, 63, 63, 63, 63, 64, 64, 64, 64, 64, 64, 64, 64, 65, 65, 65, 65, 65, 65, 65, 65, 66, 66, 66, 66, 66, 66, 67, 67, 67, 67, 67, 67, 68, 68, 68, 68, 69, 69, 69, 69, 69, 69, 70, 70, 70, 70, 70, 70, 70, 71, 71, 71, 71, 71, 71, 71, 71, 72, 72, 72, 72, 72, 72, 72, 72, 73, 73, 73, 73, 73, 73, 73, 73, 74, 74, 74, 74, 74, 75, 75, 75, 75, 75, 75, 75, 75, 76, 76, 76, 76, 76, 76, 77, 77, 77, 77, 77, 77, 77, 77, 78, 78, 78, 78, 78, 78, 78, 78, 79, 79, 79, 79, 79, 79, 79, 79, 80, 80, 80, 80, 80, 80, 80, 80, 81, 81, 81, 81, 81, 81, 81, 81, 82, 82, 82, 82, 82, 82, 83, 83, 83, 83, 83, 83, 83, 83, 84, 84, 84, 84, 84, 84, 84, 84, 85, 85, 85, 85, 85, 85, 85, 85, 86, 86, 86, 86, 86, 86, 86, 87, 87, 87, 87, 87, 87, 87, 88, 88, 88, 88, 88, 88, 88, 88, 89, 89, 89, 89, 89, 89, 89, 89, 90, 90, 90, 90, 90, 90, 90, 90, 91, 91, 91, 91, 91, 91, 92, 92, 92, 92, 92, 92, 92, 93, 93, 93, 94, 94, 94, 94, 94, 94, 95, 95, 95, 95, 95, 95, 95, 96, 96, 96, 96, 96, 96, 96, 96, 97, 97, 97, 97, 97, 97, 97, 97, 98, 98, 98, 98, 98, 98, 98, 98, 99, 99, 99, 99, 99, 99, 100, 100, 100, 100, 100, 100, 100, 101, 101, 101, 101, 101, 101, 102, 102, 102, 102, 102, 102, 102, 102, 103, 103, 103, 103, 103, 103, 103, 103, 104, 104, 104, 104, 104, 104, 104, 104, 105, 105, 105, 105, 105, 105, 105, 105, 106, 106, 106, 106, 106, 106, 106, 106, 107, 107, 107, 107, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 109, 109, 109, 109, 109, 109, 109, 109, 110, 110, 110, 110, 110, 110, 110, 110, 111, 111, 111, 111, 111, 111, 111, 111, 112, 112, 112, 112, 112, 112, 113, 113, 113, 113, 113, 113, 113, 113, 114, 114, 114, 114, 114, 114, 114, 114, 115, 115, 115, 115, 115, 115, 115, 115, 116, 116, 116, 116, 116, 116, 117, 117, 117, 117, 117, 117, 117, 118, 118, 118, 118, 119, 119, 119, 119, 119, 120, 120, 120, 120, 120, 120, 120, 121, 121, 121, 121, 121, 121, 121, 121, 122, 122, 122, 122, 122, 122, 122, 122, 123, 123, 123, 123, 123, 123, 123, 123, 124, 124, 124, 124, 124, 124, 124, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 129, 129, 129, 129, 129, 129, 129, 129, 130, 130, 130, 130, 130, 130, 130, 130, 131, 131, 131, 131, 131, 131, 131, 131, 132, 132, 132, 132, 132, 132, 132, 133, 133, 133, 133, 133, 133, 133, 134, 134, 134, 134, 134, 134, 134, 134, 135, 135, 135, 135, 135, 135, 135, 135, 136, 136, 136, 136, 136, 136, 136, 136, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 138, 138, 138, 139, 139, 139, 139, 139, 139, 139, 139, 140, 140, 140, 140, 140, 140, 140, 140, 141, 141, 141, 141, 141, 141, 142, 142, 142, 142, 142, 142, 142, 143, 143, 143, 143, 143, 144, 144, 144, 144, 145, 145, 145, 145, 145, 145, 145, 146, 146, 146, 146, 146, 146, 146, 146, 147, 147, 147, 147, 147, 147, 147, 147, 148, 148, 148, 148, 148, 148, 148, 148, 149, 149, 149, 149, 149, 149, 149, 149, 150, 150, 150, 150, 150, 151, 151, 151, 151, 151, 151, 151, 152, 152, 152, 152, 152, 152, 152, 153, 153, 153, 153, 153, 153, 153, 153, 154, 154, 154, 154, 154, 154, 154, 154, 155, 155, 155, 155, 155, 155, 155, 155, 156, 156, 156, 156, 156, 156, 156, 156, 157, 157, 157, 157, 157, 157, 157, 158, 158, 158, 158, 158, 158, 158, 159, 159, 159, 159, 159, 159, 159, 159, 160, 160, 160, 160, 160, 160, 160, 160, 161, 161, 161, 161, 161, 161, 161, 161, 162, 162, 162, 162, 162, 162, 163, 163, 163, 163, 163, 163, 163, 163, 164, 164, 164, 164, 164, 164, 164, 164, 165, 165, 165, 165, 165, 165, 165, 165, 166, 166, 166, 166, 166, 166, 166, 167, 167, 167, 167, 167, 167, 167, 168, 168, 168, 168, 169, 169, 169, 169, 169, 170, 170, 170, 170, 170, 170, 171, 171, 171, 171, 171, 171, 171, 171, 172, 172, 172, 172, 172, 172, 172, 172, 173, 173, 173, 173, 173, 173, 173, 173, 174, 174, 174, 174, 174, 174, 174, 174, 175, 175, 175, 175, 175, 176, 176, 176, 176, 176, 176, 176, 177, 177, 177, 177, 177, 177, 177, 178, 178, 178, 178, 178, 178, 178, 178, 179, 179, 179, 179, 179, 179, 179, 179, 180, 180, 180, 180, 180, 180, 180, 180, 181, 181, 181, 181, 181, 181, 181, 181, 182, 182, 182, 182, 182, 182, 182, 183, 183, 183, 183, 183, 183, 183, 184, 184, 184, 184, 184, 184, 184, 184, 185, 185, 185, 185, 185, 185, 185, 185, 186, 186, 186, 186, 186, 186, 186, 186, 187, 187, 187, 187, 187, 187, 188, 188, 188, 188, 188, 188, 188, 188, 189, 189, 189, 189, 189, 189, 189, 189, 190, 190, 190, 190, 190, 190, 190, 190, 191, 191, 191, 191, 191, 191, 191, 192, 192, 192, 192, 192, 192, 192, 193, 193, 193, 193, 194, 194, 194, 194, 194, 195, 195, 195, 195, 195, 196, 196, 196, 196, 196, 196, 196, 196, 197, 197, 197, 197, 197, 197, 197, 197, 198, 198, 198, 198, 198, 198, 198, 198, 199, 199, 199, 199, 199, 199, 199, 199, 200, 200, 200, 200, 200, 201, 201, 201, 201, 201, 201, 201, 201, 202, 202, 202, 202, 202, 202, 203, 203, 203, 203, 203, 203, 203, 203, 204, 204, 204, 204, 204, 204, 204, 204, 205, 205, 205, 205, 205, 205, 205, 205, 206, 206, 206, 206, 206, 206, 206, 206, 207, 207, 207, 207, 207, 207, 207, 207, 208, 208, 208, 208, 208, 208, 208, 208, 209, 209, 209, 209, 209, 209, 209, 209, 210, 210, 210, 210, 210, 210, 210, 210, 211, 211, 211, 211, 211, 211, 211, 211, 212, 212, 212, 212, 212, 212, 212, 212, 213, 213, 213, 213, 213, 213, 213, 213, 214, 214, 214, 214, 214, 214, 215, 215, 215, 215, 215, 215, 215, 215, 216, 216, 216, 216, 216, 217, 217, 217, 217, 217, 217, 218, 218, 218, 218, 218, 218, 218, 219, 219, 219, 219, 219, 219, 220, 220, 220, 220, 221, 221, 221, 221, 221, 221, 221, 222, 222, 222, 222, 222, 222, 222, 223, 223, 223, 223, 223, 223, 223, 223, 224, 224, 224, 224, 224, 224, 224, 225, 225, 225, 225, 226, 226, 226, 226, 226, 226, 226, 227, 227, 227, 227, 227, 227, 227, 227, 228, 228, 228, 228, 228, 228, 228, 228, 229, 229, 229, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 231, 231, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 232, 232, 233, 233, 233, 233, 233, 233, 234, 234, 234, 234, 234, 234, 234, 234, 235, 235, 235, 235, 235, 235, 235, 236, 236, 236, 236, 236, 236, 236, 237, 237, 237, 237, 237, 237, 237, 238, 238, 238, 238, 238, 238, 238, 239, 239, 239, 239, 239, 239, 239, 239, 240, 240, 240, 240, 240, 240, 240, 240, 241, 241, 241, 241, 241, 241, 241, 241, 242, 242, 242, 242, 243, 243, 243, 243, 243, 243, 244, 244, 244, 244, 244, 244, 244, 244, 245, 245, 245, 245, 245, 245, 245, 245, 246, 246, 246, 246, 246, 246, 247, 247, 247, 247, 247, 247, 247, 247, 248, 248, 248, 248, 248, 248, 248, 248, 249, 249, 249, 249, 249, 249, 249, 249, 250, 250, 250, 250, 250, 250, 250, 251, 251, 251, 251, 251, 251, 251, 252, 252, 252, 252, 252, 252, 252, 252, 253, 253, 253, 253, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 256, 256, 256, 257, 257, 257, 257, 257, 258, 258, 258, 259, 259, 259, 259, 259, 260, 260, 261, 261, 261, 261, 261, 261, 262, 262, 262, 262, 263, 263, 263, 263, 264, 264, 264, 264, 264, 265, 265, 265, 266, 266, 266, 266, 266, 266, 266, 267, 267, 267, 267, 267, 268, 268, 269, 269, 269, 269, 269, 269, 270, 270, 270, 270, 270, 271, 271, 271, 271, 271, 272, 272, 272, 272, 272, 272, 272, 273, 273, 273, 273, 273, 273, 273, 274, 274, 274, 274, 274, 274, 274, 274, 275, 275, 275, 275, 275, 275, 275, 276, 277, 277, 277, 277, 278, 278, 278, 278, 278, 278, 278, 279, 279, 279, 279, 279, 279, 279, 279, 280, 280, 280, 280, 280, 280, 280, 280, 281, 281, 281, 281, 281, 281, 281, 281, 282, 283, 283, 283, 284, 284, 284, 285, 285, 285, 285, 285, 286, 286, 286, 287, 287, 287, 287, 287, 288, 288, 288, 288, 288, 289, 289, 289, 290, 290, 290, 290, 290, 290, 290, 290, 291, 291, 291, 291, 291, 292, 292, 293, 293, 293, 293, 293, 293, 293, 294, 294, 294, 294, 294, 294, 295, 295, 295, 295, 295, 295, 295, 296, 296, 296, 296, 296, 296, 297, 297, 298, 298, 298, 298, 298, 298, 298, 299, 299, 299, 299, 299, 299, 299, 299, 300, 300, 300, 300, 300, 300, 300, 300, 301, 301, 301, 301, 301, 301, 301, 301, 302, 302, 302, 302, 302, 302, 302, 302, 303, 303, 303, 303, 303, 303, 303, 303, 304, 304, 304, 304, 304, 304, 304, 304, 305, 305, 305, 305, 305, 305, 306, 306, 306, 306, 306, 306, 306, 306, 307, 307, 307, 307, 307, 308, 308, 308, 308, 308, 308, 309, 309, 309, 309, 309, 309, 309, 310, 310, 310, 310, 310, 310, 311, 311, 311, 311, 311, 312, 312, 312, 312, 312, 312, 312, 313, 313, 313, 313, 313, 313, 313, 314, 314, 314, 314, 314, 314, 314, 314, 315, 315, 315, 315, 315, 315, 316, 316, 316, 316, 317, 317, 317, 317, 317, 317, 317, 317, 318, 318, 318, 318, 318, 318, 318, 318, 319, 319, 319, 319, 319, 319, 319, 319, 320, 320, 320, 320, 320, 320, 321, 321, 321, 321, 321, 321, 321, 321, 322, 322, 322, 322, 322, 322, 322, 322, 323, 323, 323, 323, 323, 323, 323, 323, 324, 324, 324, 324, 324, 324, 325, 325, 325, 325, 325, 325, 325, 325, 326, 326, 326, 326, 326, 326, 327, 327, 327, 327, 327, 327, 327, 327, 328, 328, 328, 328, 328, 328, 328, 329, 329, 329, 329, 329, 329, 329, 330, 330, 330, 330, 330, 330, 330, 330, 331, 331, 331, 331, 331, 331, 331, 331, 332, 332, 332, 332, 332, 332, 332, 332, 333, 333, 333, 333, 334, 334, 334, 334, 334, 334, 335, 335, 335, 335, 335, 335, 335, 335, 336, 336, 336, 336, 336, 336, 336, 336, 337, 337, 337, 337, 337, 337, 338, 338, 338, 338, 338, 338, 338, 338, 339, 339, 339, 339, 339, 339, 339, 339, 340, 340, 340, 340, 340, 340, 340, 340, 341, 341, 341, 341, 341, 341, 341, 342, 342, 342, 342, 342, 342, 342, 343, 343, 343, 343, 343, 343, 343, 343, 344, 344, 344, 344, 345, 345, 345, 345, 345, 345, 345, 346, 346, 346, 346, 347, 347, 347, 347, 348, 348, 348, 348, 349, 349, 349, 350, 350, 350, 350, 350, 350, 351, 352, 352, 352, 352, 352, 352, 352, 353, 353, 353, 354, 354, 354, 354, 354, 355, 355, 355, 355, 356, 356, 356, 356, 357, 357, 357, 357, 357, 357, 357, 358, 358, 358, 358, 359, 359, 359, 360, 360, 360, 360, 360, 360, 361, 361, 361, 361, 362, 362, 362, 362, 362, 362, 363, 363, 363, 363, 363, 363, 363, 364, 364, 364, 364, 364, 364, 364, 365, 365, 365, 365, 365, 365, 365, 366, 366, 366, 366, 366, 366, 366, 366, 368, 368, 368, 368, 368, 369, 369, 369, 369, 369, 369, 369, 370, 370, 370, 370, 370, 370, 370, 370, 371, 371, 371, 371, 371, 371, 371, 371, 372, 372, 372, 372, 372, 372, 372, 372, 374, 374, 374, 375, 375, 375, 376, 376, 376, 376, 376, 376, 376, 377, 377, 378, 378, 378, 378, 378, 379, 379, 379, 379, 380, 380, 380, 380, 381, 381, 381, 381, 381, 381, 382, 382, 382, 382, 382, 383, 383, 383, 383, 384, 384, 384, 384, 384, 384, 384, 385, 385, 385, 385, 385, 385, 386, 386, 387, 387, 387, 387, 387, 387, 387, 387, 388, 388, 388, 388, 388, 388, 389, 390, 390, 390, 390, 390, 390, 390, 390, 391, 391, 391, 391, 391, 391, 391, 391, 392, 392, 392, 392, 392, 392, 392, 392, 393, 393, 393, 393, 393, 393, 393, 393, 394, 394, 394, 394, 394, 394, 394, 394, 395, 395, 395, 395, 395, 395, 395, 395, 396, 396, 396, 396, 396, 396, 396, 397, 397, 397, 397, 397, 397, 397, 398, 398, 398, 398, 398, 398, 398, 398, 399, 399, 399, 399, 399, 400, 400, 400, 400, 400, 400, 401, 401, 401, 401, 401, 401, 402, 402, 402, 402, 402, 403, 403, 403, 403, 403, 403, 403, 404, 404, 404, 404, 404, 404, 404, 405, 405, 405, 405, 405, 405, 405, 406, 406, 406, 406, 406, 406, 406, 406, 407, 407, 407, 407, 407, 408, 408, 408, 408, 408, 409, 409, 409, 409, 409, 409, 409, 409, 410, 410, 410, 410, 410, 410, 410, 410, 411, 411, 411, 411, 411, 411, 411, 412, 412, 412, 412, 412, 412, 412, 413, 413, 413, 413, 413, 413, 413, 413, 414, 414, 414, 414, 414, 414, 414, 414, 415, 415, 415, 415, 415, 415, 415, 415, 416, 416, 416, 416, 416, 416, 417, 417, 417, 417, 417, 417, 417, 417, 418, 418, 418, 418, 418, 418, 419, 419, 419, 419, 419, 419, 419, 420, 420, 420, 420, 420, 420, 420, 421, 421, 421, 421, 421, 421, 421, 421, 422, 422, 422, 422, 422, 422, 422, 422, 423, 423, 423, 423, 423, 423, 423, 423, 424, 424, 424, 424, 424, 424, 425, 425, 425, 425, 426, 426, 426, 426, 426, 426, 426, 426, 427, 427, 427, 427, 427, 427, 427, 427, 428, 428, 428, 428, 428, 428, 428, 428, 429, 429, 429, 429, 429, 429, 430, 430, 430, 430, 430, 430, 430, 430, 431, 431, 431, 431, 431, 431, 431, 431, 432, 432, 432, 432, 432, 432, 432, 432, 433, 433, 433, 433, 433, 433, 434, 434, 434, 434, 434, 434, 434, 434, 435, 435, 435, 435, 435, 435, 436, 436, 436, 436, 436, 437, 437, 437, 437, 437, 437, 437, 437, 438, 438, 438, 439, 439, 439, 439, 440, 440, 440, 440, 441, 441, 441, 441, 442, 442, 442, 442, 443, 443, 444, 444, 444, 444, 444, 444, 444, 444, 445, 445, 446, 446, 446, 446, 446, 447, 447, 447, 447, 448, 448, 448, 448, 448, 449, 449, 449, 449, 449, 449, 449, 450, 450, 451, 451, 451, 451, 451, 452, 452, 452, 452, 453, 453, 453, 453, 454, 454, 454, 454, 454, 454, 454, 454, 455, 455, 455, 455, 455, 455, 456, 456, 456, 456, 456, 456, 456, 456, 457, 457, 457, 457, 457, 457, 457, 458, 458, 458, 458, 458, 458, 459, 460, 460, 460, 460, 460, 460, 461, 461, 461, 461, 461, 461, 461, 462, 462, 462, 462, 462, 462, 462, 462, 463, 463, 463, 463, 463, 463, 463, 463, 464, 464, 464, 464, 464, 464, 465, 466, 466, 466, 466, 467, 467, 468, 468, 468, 468, 468, 468, 468, 469, 469, 469, 470, 470, 470, 470, 471, 471, 471, 471, 472, 472, 472, 472, 473, 473, 473, 473, 473, 473, 474, 474, 474, 474, 474, 475, 475, 475, 475, 475, 476, 476, 476, 476, 476, 476, 477, 477, 477, 477, 477, 478, 478, 478, 478, 479, 479, 479, 479, 479, 479, 479, 479, 480, 480, 480, 480, 481, 481, 481, 482, 482, 482, 482, 482, 482, 482, 482, 483, 483, 483, 483, 483, 483, 483, 483, 484, 484, 484, 484, 484, 484, 484, 484, 485, 485, 485, 485, 485, 485, 485, 485, 486, 486, 486, 486, 486, 486, 486, 486, 487, 487, 487, 487, 487, 487, 487, 487, 488, 488, 488, 488, 488, 488, 489, 489, 489, 489, 489, 489, 489, 489, 490, 490, 490, 490, 490, 490, 491, 491, 491, 491, 491, 491, 492, 492, 492, 492, 492, 492, 492, 493, 493, 493, 493, 493, 493, 494, 494, 494, 494, 495, 495, 495, 495, 495, 495, 495, 496, 496, 496, 496, 496, 496, 496, 496, 497, 497, 497, 497, 497, 497, 497, 498, 498, 498, 498, 498, 498, 498, 498, 499, 499, 499, 499, 499, 500, 500, 500, 500, 500, 501, 501, 501, 501, 501, 501, 501, 501, 502, 502, 502, 502, 502, 502, 502, 502, 503, 503, 503, 503, 503, 503, 504, 504, 504, 504, 504, 504, 504, 504, 505, 505, 505, 505, 505, 505, 505, 505, 506, 506, 506, 506, 506, 506, 506, 506, 507, 507, 507, 507, 507, 507, 507, 508, 508, 508, 508, 508, 508, 508, 509, 509, 509, 509, 509, 509, 509, 509, 510, 510, 510, 510, 510, 510, 511, 511, 511, 511, 511, 511, 511, 512, 512, 512, 512, 512, 512, 512, 513, 513, 513, 513, 513, 513, 513, 513, 514, 514, 514, 514, 514, 514, 514, 514, 515, 515, 515, 515, 515, 515, 515, 515, 516, 516, 516, 516, 516, 517, 517, 517, 517, 517, 518, 518, 518, 518, 518, 518, 518, 518, 519, 519, 519, 519, 519, 519, 519, 519, 520, 520, 520, 520, 520, 520, 520, 521, 521, 521, 521, 521, 521, 521, 522, 522, 522, 522, 522, 522, 522, 522, 523, 523, 523, 523, 523, 523, 523, 523, 524, 524, 524, 524, 524, 524, 524, 524, 525, 525, 525, 525, 525, 525, 526, 526, 526, 526, 526, 526, 526, 526, 527, 527, 527, 527, 527, 528, 528, 528, 528, 528, 528, 529, 529, 529, 529, 529, 529, 529, 530, 530, 530, 531, 531, 531, 531, 531, 532, 532, 533, 533, 533, 533, 533, 533, 534, 534, 535, 535, 535, 535, 536, 536, 536, 536, 536, 536, 536, 537, 538, 538, 538, 538, 538, 539, 539, 539, 539, 540, 540, 540, 540, 540, 540, 541, 541, 541, 541, 541, 541, 541, 541, 542, 543, 543, 543, 543, 544, 544, 544, 544, 544, 544, 545, 545, 545, 545, 546, 546, 546, 546, 546, 546, 546, 547, 547, 547, 547, 547, 547, 547, 548, 548, 548, 548, 548, 548, 548, 548, 549, 549, 549, 549, 549, 549, 549, 550, 550, 550, 550, 551, 552, 552, 552, 552, 552, 552, 552, 552, 553, 553, 553, 553, 553, 553, 553, 554, 554, 554, 554, 554, 554, 554, 554, 555, 555, 555, 555, 555, 555, 555, 555, 556, 556, 556, 556, 557, 558, 558, 558, 558, 559, 559, 559, 559, 560, 560, 560, 560, 560, 561, 561, 561, 562, 562, 562, 562, 562, 563, 563, 563, 564, 564, 564, 564, 564, 564, 565, 565, 565, 565, 565, 566, 566, 566, 566, 567, 567, 567, 567, 567, 567, 567, 568, 568, 568, 568, 568, 569, 569, 569, 569, 570, 570, 570, 570, 570, 570, 571, 571, 571, 571, 571, 571, 571, 571, 572, 572, 573, 573, 573, 573, 573, 574, 574, 574, 574, 574, 574, 574, 574, 575, 575, 575, 575, 575, 575, 575, 575, 576, 576, 576, 576, 576, 576, 576, 576, 577, 577, 577, 577, 577, 577, 577, 577, 578, 578, 578, 578, 578, 578, 578, 578, 579, 579, 579, 579, 579, 579, 579, 579, 580, 580, 580, 580, 580, 580, 581, 581, 581, 581, 581, 581, 581, 581, 582, 582, 582, 582, 582, 582, 583, 583, 583, 583, 583, 583, 584, 584, 584, 584, 584, 584, 584, 585, 585, 585, 585, 585, 585, 586, 586, 586, 586, 587, 587, 587, 587, 587, 587, 587, 588, 588, 588, 588, 588, 588, 588, 589, 589, 589, 589, 589, 589, 589, 589, 590, 590, 590, 590, 590, 590, 590, 590, 591, 591, 591, 591, 592, 592, 592, 592, 592, 592, 593, 593, 593, 593, 593, 593, 593, 593, 594, 594, 594, 594, 594, 594, 594, 594, 595, 595, 595, 595, 595, 595, 596, 596, 596, 596, 596, 596, 596, 596, 597, 597, 597, 597, 597, 597, 597, 597, 598, 598, 598, 598, 598, 598, 598, 598, 599, 599, 599, 599, 599, 599, 599, 600, 600, 600, 600, 600, 600, 600, 601, 601, 601, 601, 601, 601, 601, 601, 602, 602, 602, 602, 602, 602, 603, 603, 603, 603, 603, 603, 603, 604, 604, 604, 604, 604, 604, 604, 605, 605, 605, 605, 605, 605, 605, 605, 606, 606, 606, 606, 606, 606, 606, 606, 607, 607, 607, 607, 607, 607, 607, 607, 608, 608, 608, 608, 608, 609, 609, 609, 609, 609, 610, 610, 610, 610, 610, 610, 610, 610, 611, 611, 611, 611, 611, 611, 611, 611, 612, 612, 612, 612, 612, 612, 613, 613, 613, 613, 613, 613, 613, 613, 614, 614, 614, 614, 614, 614, 614, 614, 615, 615, 615, 615, 615, 615, 615, 615, 616, 616, 616, 616, 616, 616, 616, 617, 617, 617, 617, 617, 617, 617, 618, 618, 618, 618, 618, 618, 618, 618, 619, 619, 619, 619, 620, 620, 620, 620, 620, 620, 620, 621, 621, 621, 621, 621, 622, 622, 622, 622, 623, 623, 623, 623, 623, 624, 624, 625, 625, 625, 625, 625, 626, 626, 626, 627, 627, 627, 627, 627, 628, 628, 628, 628, 628, 629, 629, 629, 630, 630, 630, 630, 630, 631, 631, 631, 632, 632, 632, 632, 632, 632, 632, 633, 633, 633, 633, 633, 633, 634, 635, 635, 635, 635, 635, 635, 636, 636, 636, 636, 636, 637, 637, 637, 637, 637, 638, 638, 638, 638, 638, 638, 638, 639, 639, 639, 639, 639, 639, 639, 640, 640, 640, 640, 640, 640, 640, 640, 641, 641, 641, 641, 641, 641, 641, 642, 642, 643, 643, 643, 644, 644, 644, 644, 644, 644, 644, 645, 645, 645, 645, 645, 645, 645, 645, 646, 646, 646, 646, 646, 646, 646, 646, 647, 647, 647, 647, 647, 647, 647, 647, 648, 648, 649, 649, 649, 650, 650, 650, 651, 651, 651, 651, 651, 652, 652, 652, 652, 653, 653, 653, 653, 654, 654, 654, 654, 655, 655, 655, 656, 656, 656, 656, 656, 656, 657, 657, 657, 657, 657, 657, 658, 658, 658, 659, 659, 659, 659, 659, 659, 659, 659, 660, 660, 660, 660, 660, 661, 661, 661, 662, 662, 662, 662, 662, 662, 662, 663, 663, 663, 663, 663, 663, 664, 664, 665, 665, 665, 665, 665, 665, 665, 666, 666, 666, 666, 666, 666, 666, 666, 667, 667, 667, 667, 667, 667, 667, 667, 668, 668, 668, 668, 668, 668, 668, 668, 669, 669, 669, 669, 669, 669, 669, 669, 670, 670, 670, 670, 670, 670, 670, 670, 671, 671, 671, 671, 671, 671, 671, 671, 672, 672, 672, 672, 672, 672, 673, 673, 673, 673, 673, 673, 673, 673, 674, 674, 674, 674, 674, 675, 675, 675, 675, 675, 675, 676, 676, 676, 676, 676, 676, 676, 677, 677, 677, 677, 677, 677, 678, 678, 678, 678, 678, 679, 679, 679, 679, 679, 679, 679, 680, 680, 680, 680, 680, 680, 680, 681, 681, 681, 681, 681, 681, 681, 681, 682, 682, 682, 682, 682, 682, 683, 683, 683, 683, 684, 684, 684, 684, 684, 684, 684, 684, 685, 685, 685, 685, 685, 685, 685, 685, 686, 686, 686, 686, 686, 686, 686, 686, 687, 687, 687, 687, 687, 687, 688, 688, 688, 688, 688, 688, 688, 688, 689, 689, 689, 689, 689, 689, 689, 689, 690, 690, 690, 690, 690, 690, 690, 690, 691, 691, 691, 691, 691, 691, 692, 692, 692, 692, 692, 692, 692, 692, 693, 693, 693, 693, 693, 693, 694, 694, 694, 694, 694, 694, 694, 694, 695, 695, 695, 695, 695, 695, 695, 696, 696, 696, 696, 696, 696, 696, 697, 697, 697, 697, 697, 697, 697, 697, 698, 698, 698, 698, 698, 698, 698, 698, 699, 699, 699, 699, 699, 699, 699, 699, 700, 700, 700, 700, 701, 701, 701, 701, 701, 701, 702, 702, 702, 702, 702, 702, 702, 702, 703, 703, 703, 703, 703, 703, 703, 703, 704, 704, 704, 704, 704, 704, 705, 705, 705, 705, 705, 705, 705, 705, 706, 706, 706, 706, 706, 706, 706, 706, 707, 707, 707, 707, 707, 707, 707, 707, 708, 708, 708, 708, 708, 708, 708, 709, 709, 709, 709, 709, 709, 709, 710, 710, 710, 710, 710, 710, 710, 710, 711, 711, 711, 711, 712, 712, 712, 712, 712, 712, 712, 713, 713, 713, 713, 714, 714, 714, 714, 715, 715, 715, 715, 716, 716, 716, 717, 717, 717, 717, 717, 717, 718, 719, 719, 719, 719, 719, 719, 719, 720, 720, 720, 721, 721, 721, 721, 721, 722, 722, 722, 722, 723, 723, 723, 723, 724, 724, 724, 724, 724, 724, 724, 725, 725, 725, 725, 726, 726, 726, 727, 727, 727, 727, 727, 727, 728, 728, 728, 728, 729, 729, 729, 729, 729, 729, 730, 730, 730, 730, 730, 730, 730, 731, 731, 731, 731, 731, 731, 731, 732, 732, 732, 732, 732, 732, 732, 733, 733, 733, 733, 733, 733, 733, 733, 735, 735, 735, 735, 735, 736, 736, 736, 736, 736, 736, 736, 737, 737, 737, 737, 737, 737, 737, 737, 738, 738, 738, 738, 738, 738, 738, 738, 739, 739, 739, 739, 739, 739, 739, 739, 741, 741, 741, 742, 742, 742, 743, 743, 743, 743, 743, 743, 743, 744, 744, 745, 745, 745, 745, 745, 746, 746, 746, 746, 747, 747, 747, 747, 748, 748, 748, 748, 748, 748, 749, 749, 749, 749, 749, 750, 750, 750, 750, 751, 751, 751, 751, 751, 751, 751, 752, 752, 752, 752, 752, 752, 753, 753, 754, 754, 754, 754, 754, 754, 754, 754, 755, 755, 755, 755, 755, 755, 756, 757, 757, 757, 757, 757, 757, 757, 757, 758, 758, 758, 758, 758, 758, 758, 758, 759, 759, 759, 759, 759, 759, 759, 759, 760, 760, 760, 760, 760, 760, 760, 760, 761, 761, 761, 761, 761, 761, 761, 761, 762, 762, 762, 762, 762, 762, 762, 762, 763, 763, 763, 763, 763, 763, 763, 764, 764, 764, 764, 764, 764, 764, 765, 765, 765, 765, 765, 765, 765, 765, 766, 766, 766, 766, 766, 767, 767, 767, 767, 767, 767, 768, 768, 768, 768, 768, 768, 769, 769, 769, 769, 769, 770, 770, 770, 770, 770, 770, 770, 771, 771, 771, 771, 771, 771, 771, 772, 772, 772, 772, 772, 772, 772, 773, 773, 773, 773, 773, 773, 773, 773, 774, 774, 774, 774, 774, 775, 775, 775, 775, 775, 776, 776, 776, 776, 776, 776, 776, 776, 777, 777, 777, 777, 777, 777, 777, 777, 778, 778, 778, 778, 778, 778, 778, 779, 779, 779, 779, 779, 779, 779, 780, 780, 780, 780, 780, 780, 780, 780, 781, 781, 781, 781, 781, 781, 781, 781, 782, 782, 782, 782, 782, 782, 782, 782, 783, 783, 783, 783, 783, 783, 784, 784, 784, 784, 784, 784, 784, 784, 785, 785, 785, 785, 785, 785, 786, 786, 786, 786, 786, 786, 786, 787, 787, 787, 787, 787, 787, 787, 788, 788, 788, 788, 788, 788, 788, 788, 789, 789, 789, 789, 789, 789, 789, 789, 790, 790, 790, 790, 790, 790, 790, 790, 791, 791, 791, 791, 791, 791, 792, 792, 792, 792, 793, 793, 793, 793, 793, 793, 793, 793, 794, 794, 794, 794, 794, 794, 794, 794, 795, 795, 795, 795, 795, 795, 795, 795, 796, 796, 796, 796, 796, 796, 797, 797, 797, 797, 797, 797, 797, 797, 798, 798, 798, 798, 798, 798, 798, 798, 799, 799, 799, 799, 799, 799, 799, 799, 800, 800, 800, 800, 800, 800, 801, 801, 801, 801, 801, 801, 801, 801, 802, 802, 802, 802, 802, 802, 803, 803, 803, 803, 803, 804, 804, 804, 804, 804, 804, 804, 804, 805, 805, 805, 806, 806, 806, 806, 807, 807, 807, 807, 808, 808, 808, 808, 809, 809, 809, 809, 810, 810, 811, 811, 811, 811, 811, 811, 811, 811, 812, 812, 813, 813, 813, 813, 813, 814, 814, 814, 814, 815, 815, 815, 815, 815, 816, 816, 816, 816, 816, 816, 816, 817, 817, 818, 818, 818, 818, 818, 819, 819, 819, 819, 820, 820, 820, 820, 821, 821, 821, 821, 821, 821, 821, 821, 822, 822, 822, 822, 822, 822, 823, 823, 823, 823, 823, 823, 823, 823, 824, 824, 824, 824, 824, 824, 824, 825, 825, 825, 825, 825, 825, 826, 827, 827, 827, 827, 827, 827, 828, 828, 828, 828, 828, 828, 828, 829, 829, 829, 829, 829, 829, 829, 829, 830, 830, 830, 830, 830, 830, 830, 830, 831, 831, 831, 831, 831, 831, 832, 833, 833, 833, 833, 834, 834, 835, 835, 835, 835, 835, 835, 835, 836, 836, 836, 837, 837, 837, 837, 838, 838, 838, 838, 839, 839, 839, 839, 840, 840, 840, 840, 840, 840, 841, 841, 841, 841, 841, 842, 842, 842, 842, 842, 843, 843, 843, 843, 843, 843, 844, 844, 844, 844, 844, 845, 845, 845, 845, 846, 846, 846, 846, 846, 846, 846, 846, 847, 847, 847, 847, 848, 848, 848, 849, 849, 849, 849, 849, 849, 849, 849, 850, 850, 850, 850, 850, 850, 850, 850, 851, 851, 851, 851, 851, 851, 851, 851, 852, 852, 852, 852, 852, 852, 857, 857, 857, 857, 857, 858, 858, 858, 858, 858, 858, 858, 858, 859, 859, 859, 859, 859, 860, 860, 860, 860, 860, 861, 861, 861, 861, 861, 861, 861, 861, 862, 862, 862, 862, 862, 862, 862, 862, 863, 863, 863, 863, 863, 863, 863, 864, 864, 864, 864, 864, 864, 864, 865, 865, 865, 865, 865, 865, 865, 865, 866, 866, 866, 866, 866, 866, 866, 866, 867, 867, 867, 867, 867, 867, 867, 867, 868, 868, 868, 868, 868, 868, 869, 869, 869, 869, 869, 869, 869, 869, 870, 870, 870, 870, 870, 870, 871, 871, 871, 871, 871, 871, 871, 872, 872, 872, 872, 872, 872, 872, 873, 873, 873, 873, 873, 873, 873, 873, 874, 874, 874, 874, 874, 874, 874, 874, 875, 875, 875, 875, 875, 875, 875, 875, 876, 876, 876, 876, 876, 876, 877, 877, 877, 877, 878, 878, 878, 878, 878, 878, 878, 878, 879, 879, 879, 879, 879, 879, 879, 879, 880, 880, 880, 880, 880, 880, 880, 880, 881, 881, 881, 881, 881, 881, 882, 882, 882, 882, 882, 882, 882, 882, 883, 883, 883, 883, 883, 883, 883, 883, 884, 884, 884, 884, 884, 884, 884, 884, 885, 885, 885, 885, 885, 885, 886, 886, 886, 886, 886, 886, 886, 886, 887, 887, 887, 887, 887, 887, 888, 888, 888, 888, 888, 889, 889, 889, 889, 889, 889, 889, 889, 890, 890, 890, 891, 891, 891, 891, 892, 892, 892, 892, 893, 893, 893, 893, 894, 894, 894, 894, 895, 895, 895, 895, 895, 896, 896, 896, 896, 896, 896, 897, 897, 898, 898, 898, 898, 899, 899, 899, 900, 900, 900, 901, 901, 901, 901, 901, 901, 902, 902, 902, 902, 902, 902, 903, 903, 904, 904, 904, 904, 904, 904, 905, 905, 905, 905, 906, 906, 906, 906, 906, 906, 907, 907, 907, 907, 907, 907, 907, 908, 908, 908, 908, 908, 908, 908, 909, 909, 909, 909, 909, 909, 909, 909, 910, 910, 910, 910, 910, 910, 910, 910, 911, 911, 911, 911, 911, 911, 911, 911, 912, 912, 912, 912, 912, 912, 912, 912, 913, 913, 913, 913, 913, 913, 913, 914, 914, 914, 914, 914, 914, 915, 915, 915, 915, 915, 915, 915, 916, 916, 916, 916, 916, 916, 916, 917, 917, 917, 917, 917, 917, 917, 917, 919, 919, 919, 919, 919, 919, 920, 920, 920, 920, 920, 920, 921, 921, 921, 921, 921, 921, 921, 921, 922, 922, 922, 922, 922, 922, 922, 922, 923, 923, 923, 923, 923, 923, 923, 923, 925, 925, 925, 925, 925, 926, 926, 926, 926, 927, 927, 927, 927, 927, 928, 928, 928, 929, 929, 929, 929, 929, 929, 930, 930, 930, 930, 930, 931, 931, 931, 931, 931, 932, 932, 932, 932, 933, 933, 933, 933, 934, 934, 934, 934, 934, 935, 935, 935, 935, 935, 935, 936, 936, 936, 936, 937, 937, 937, 937, 937, 937, 937, 938, 938, 938, 938, 938, 938, 938, 938, 939, 939, 940, 940, 940, 940, 940, 940, 940, 940, 941, 941, 941, 941, 941, 941, 941, 942};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 1561;
localparam integer sub_instructions = 6;
localparam longint Inst[0:1560][0:5] = '{{64'h0, 64'h0, 64'hb4c0000000000000, 64'h2963c0780002c8, 64'he0d3b9a34e870a58, 64'h10190a4069},{64'h58170000d5bc0, 64'h149a90e64a00024, 64'h69c0000000000000, 64'hba574b95d77aff61, 64'h30a613a75f4e9d8e, 64'hd40007615},{64'h13000000000, 64'hf6a2ec5ca20000, 64'h0, 64'h4b69a7012f14b4bc, 64'h18b0f162c3c5d85, 64'h0},{64'h130000, 64'hf6b9958da80048, 64'h0, 64'h406cbdd8603274, 64'h58d3800000000d38, 64'hcb13b75f6},{64'h1300000000000000, 64'h9b2d1065640000, 64'h0, 64'hf88003e2, 64'h1d8e034be50d2f8, 64'h1018002860},{64'h0, 64'h16a3d4d441c0000, 64'h0, 64'h1e0000000001e0, 64'hca39431be0006f8, 64'h28e5},{64'h0, 64'h1075a4d5b140000, 64'h6780000000000000, 64'h32c000cb000344, 64'ha4000290000000, 64'hd199f0000},{64'h0, 64'h9ba2d493980000, 64'h0, 64'h49a0012f00033c, 64'h9000000000001268, 64'hd225f33e6},{64'h0, 64'h128268b42ac0000, 64'h0, 64'h3fc000ff000000, 64'h815d8003e4000f90, 64'h700005763},{64'h0, 64'hb4525073140000, 64'h7fc0000000000000, 64'h3f4000fd1ff3f4, 64'h760001d8000000, 64'h0},{64'h0, 64'he65eb695240000, 64'h0, 64'he800000000000000, 64'h7424e1da3a0768, 64'h49c0},{64'h0, 64'hd5458f641c0000, 64'h0, 64'h542a80015d000000, 64'h1548002a8aa55d1, 64'h0},{64'h0, 64'hf649d175200000, 64'h0, 64'h564ac0000000062c, 64'h4b49592d2, 64'h18b8000000},{64'h0, 64'h127c5f0722c0000, 64'h0, 64'h4b650ca1800000, 64'hd80003600012d8, 64'h3600},{64'h0, 64'h149b94c54a00000, 64'haa40000000000000, 64'h3a00000000000296, 64'h9d000000000a59, 64'h15530560a0},{64'h0, 64'ha4a2f165a00000, 64'h0, 64'h416, 64'h318b2b60000018b0, 64'h10600056c8},{64'h0, 64'hbb22cd54180000, 64'h0, 64'h1f200000000000, 64'h1592b7564adc7c8, 64'h5640},{64'h0, 64'h1283dae53140000, 64'h0, 64'hf934e0007c800000, 64'hd399633e000cf8, 64'hcb0000000},{64'h0, 64'hd45232641c0000, 64'h99c0000000000000, 64'h4ce001338002a8, 64'hfd800000000000, 64'haa8003f60},{64'h0, 64'hc55e54922c0000, 64'h0, 64'h60a001829f161a, 64'h406000000, 64'h1019f261c0},{64'h0, 64'hab26b493900000, 64'h3a00000000000000, 64'h1e037c74000622, 64'h1be000000, 64'h78b120000},{64'h0, 64'h1375e89b2240000, 64'h0, 64'h360000d825e61a, 64'h7c00000000000000, 64'h189b0e6269},{64'h0, 64'hbad249b2900000, 64'h0, 64'h586000000004ac, 64'h586001618, 64'h9f25727c0},{64'h0, 64'h12741c9b2900000, 64'h4e80000000000000, 64'h126999332, 64'heca5800000001268, 64'h2964},{64'h0, 64'hbbdaac55200000, 64'h0, 64'h4800000000000000, 64'he8a400041851d061, 64'h7d00028e3},{64'h0, 64'hb4458f541c0000, 64'h6980000000000000, 64'h56400159000574, 64'h2980015d0, 64'hd38002980},{64'h0, 64'h8bb95495a00000, 64'h0, 64'hf532c7d40000032c, 64'h154b1f000001549, 64'h63e0},{64'h0, 64'hd54e3065a40000, 64'h4e40000000000000, 64'h344, 64'h8cd200063e000000, 64'hd213a63e6},{64'h0, 64'h9bb10bb3940000, 64'h0, 64'h4047c901000000, 64'h8d340e33e4000000, 64'h4d03},{64'h0, 64'h137524d5b140000, 64'h7f80000000000000, 64'h3fc0000000034e, 64'ha78f029e3c0000, 64'h3500},{64'h0, 64'hf6de4e62ac0000, 64'h0, 64'hff800000, 64'h1288e04a2c39870, 64'h1000e00000},{64'h0, 64'h107b528a3980000, 64'hb0c0000000000000, 64'h5b2986a12d800298, 64'h1476305350810762, 64'h1623054088},{64'h180001c040000, 64'h7148b528bc180014, 64'h57923d9c69a8af59, 64'h297aec785ab576, 64'had638f134f4f0788, 64'hd59ac4076},{64'h60100001c000000, 64'hb09ac1ab40005000, 64'h4e533d9e4c30f8b9, 64'h575c5c788f04be, 64'he8a6558275c5c000, 64'hd44f24c04},{64'h10a00000601c0, 64'hb0bb800000000000, 64'h6f94aa6c753cb369, 64'h430c58a5e184bd, 64'h68adb161e3c5a000, 64'h1ad000330d},{64'h6000070000, 64'heab44da000004014, 64'h510a2e184c5cb891, 64'h5e2883b501e0f3e4, 64'hcc000001da978d3e, 64'h9dd4432d7},{64'h601407000000100, 64'hb117cdc000000000, 64'h80d622d25c48b7a9, 64'he128e80ca38f13e3, 64'hb501d442879392fc, 64'ha22ad49ca},{64'h638004000000140, 64'h30b4bd5798000000, 64'h52123d1066d4b889, 64'ha3000000a419f1e1, 64'h58a1d47b2e68c6fd, 64'hd000032e6},{64'h1c00000060000, 64'h1000000000004280, 64'h97d43dd4b73cb1a9, 64'h42348938cb59f49c, 64'he8cf2ba291508d21, 64'hcfda3b3ca},{64'he000000010000000, 64'h70d5b15178005018, 64'h7e5034a64b54f8b9, 64'hdf49b9687021259a, 64'h7e00000200968700, 64'h12fdfa3496},{64'h700006000050000, 64'hf09bcde000000010, 64'haa108d2a6c3898b1, 64'hf129a52cff4ec1d8, 64'hf15dcdf4267c4f95, 64'h6faa91c17},{64'h100000007014c, 64'h709bb51178000000, 64'h7eb29e2a4b2cf871, 64'h624c44e8fd4e93ff, 64'h7d5b93a1d93a55ba, 64'h750df1d23},{64'h401805380000000, 64'h5136ca3062d20000, 64'h818a33d45c54d8a9, 64'hedd54aed031382aa, 64'h69275551d1aa8744, 64'h18d1392acc},{64'h1006014070000, 64'h549aad17a0000000, 64'h95cf249a5c4cf8b1, 64'h572a96555d5954b4, 64'h352ba4d553934aa6, 64'h12d8004b09},{64'h5310000000, 64'h14f5b57598007000, 64'hc216321858b098b9, 64'h5acad6c584000362, 64'hbd5f36b57cdad2b6, 64'h18be5c4b89},{64'h60140001c040000, 64'hf0f6b997a0000000, 64'hc5493aa66c4cb659, 64'h4b7530a1e07552, 64'ha8d86ca3614ed038, 64'h18b00060ea},{64'h60000001c0, 64'h715822ebb0005010, 64'hc44f36267c289869, 64'hf056c97d5b20c297, 64'h487800062e97c9d4, 64'h15560d60bc},{64'h600007000000000, 64'hf1162ef378005010, 64'h6992352a54d49871, 64'hf41f4c7d5bb1f56e, 64'h9d5b6b31f43d18b4, 64'h1066b34196},{64'h7014c0010000000, 64'hb0bbd67178000000, 64'h65542d9c4924ed49, 64'h1f3654da1f137c, 64'hc9594fb56faca000, 64'h7d9b432e7},{64'h400007018050000, 64'h30bade6000000000, 64'hc14a261056a4d4b1, 64'h6834fc147ce683fe, 64'ha0cb6004d2800cfe, 64'h1b40004d2d},{64'h400000000060140, 64'h5cb45e6000007000, 64'h7c8db3e26ac4b851, 64'h61e39d33f0e4cf, 64'h14fdf1360cc3c738, 64'haaf1360cc},{64'h1c00000060000, 64'h24d4ce0000005010, 64'h808a5bae5c549879, 64'h1229680982d4c62c, 64'h5ca6158407c48d43, 64'hf95a861dc},{64'h300800010000140, 64'ha379aec000006380, 64'h97cd962ac0412179, 64'he1bfc995d9941d1, 64'h102ebb409c3cca0, 64'h1894f181c0},{64'he000801000050000, 64'hf115560000006190, 64'hd694682e4c3cd899, 64'hc4288d68d875a1e2, 64'h4f6214358f3c49e6, 64'h18755fcbfc},{64'h2000005190400000, 64'h3179d6600000601c, 64'h126e2cf030b161, 64'h58d87c5edc95e372, 64'h82ad9f04ec7c161d, 64'h12bd5d27d9},{64'h600400000071940, 64'hf0f6800000002010, 64'hc22685b54d871, 64'h6528e58126e18b33, 64'hd8a5d98ab7ad8f91, 64'hdfdf3277a},{64'h1825380000080, 64'h70f5800000003010, 64'h51c980246c4cd889, 64'hcb52aeca194c289, 64'h10d4b5a28f512a46, 64'h10875a1f55},{64'h140000c0601c0, 64'hf0d4dc0000004008, 64'h67cba06a5c309299, 64'h6b1c368d59547d75, 64'h48cbb6b299aa8cfb, 64'hd3d491e5b},{64'h4004061140001c0, 64'hb116a41310000000, 64'h523780d87c3cd859, 64'ha3beb001271a432d, 64'h418fe4e32f68d54d, 64'h1901502b65},{64'h4519c00000000000, 64'h30b4d40000004018, 64'h14685e6c20f851, 64'h1434938d0921d43a, 64'h82d2660e3f81471a, 64'h9d6053476},{64'h638002010050040, 64'h6c00000000003000, 64'h7e9034d257d091a9, 64'ha83e56e9014e0c25, 64'hfc71e68bf86ec805, 64'h1674ed3f87},{64'h2010c3000000142, 64'hde9080000000001c, 64'h3b2abba27c2cb899, 64'h3b1c0000a6f0e3fd, 64'hecfe6001e153f09d, 64'h187b0e3514},{64'h501c04080000080, 64'h7000000000006180, 64'hc1115e2a9434d891, 64'he9e08000761051d3, 64'hbc706704a33a7874, 64'h1004eae0c9},{64'h500007000240000, 64'hf17900000000610c, 64'h143e145c2c8da9, 64'hab5555572dcf91e2, 64'h6d82d063563e8765, 64'h1626bcaad9},{64'h6000005088000000, 64'h70b0000000004018, 64'h978fae2c5c38d169, 64'h57caf4ec790f04c0, 64'h632e13c2764e878e, 64'hd665bb579},{64'h300000000010080, 64'h30c0000000000010, 64'h9356be295c39f369, 64'h4d62eaa4d8f23363, 64'h7337ea962ec618ba, 64'h191b172759},{64'h2200c00014000000, 64'h6b36de2000000010, 64'had904c9c5c3cb841, 64'h7962d9e49dc00418, 64'h3783c0059569d062, 64'h1391b46b55},{64'h4014001800, 64'h2770000000000008, 64'h97e2d00a09889, 64'hfa1db8615b717ecc, 64'he9021ac4f06b12f4, 64'h15c36741b3},{64'h201460000000180, 64'hb0f6a6c800000010, 64'hadf158586c38b899, 64'haa298aa8a5aba407, 64'h8159ec749dacf2fa, 64'h1302aa55b9},{64'h100000000020000, 64'h160000000000000c, 64'h684dae2299ca9844, 64'h4d07c4da542284, 64'hcc7de683e2000cbe, 64'hb99a237f5},{64'h428066000000080, 64'h5337440000000000, 64'h9692686a6b20cbb9, 64'h2a4547f4fea0f4d1, 64'h315d59ec019a6a16, 64'h1260004069},{64'h100000014600000, 64'h28b4000000004008, 64'h7e95562e5c449299, 64'h4b5c3efd9fa296, 64'h34f9d5860d384fd8, 64'hfd55961f5},{64'h500006188000040, 64'h70b0800000004000, 64'h4dd0be215a36c979, 64'h12b514dd5b8e1299, 64'h8c6fd002b1384f8f, 64'h154ebc2c85},{64'h406110a30000, 64'h1579a4000000001c, 64'h8ad4361e7ab4f859, 64'hfa7598b9362b577, 64'hc89c9504c1b115bf, 64'h1621501bf3},{64'hc000180, 64'hd4ac2000004094, 64'h93cf40984c54d700, 64'h12589c48a24df40d, 64'hf0de0004dc37d27b, 64'h9ccf2e356},{64'h50100000c060040, 64'h9957ce2000000008, 64'hb2102de04c38b859, 64'h4eddb0cad47373, 64'hc926df349bdb12f8, 64'haeec92bf9},{64'h10a0000021980, 64'hd006a000000000, 64'h530b861e49dca900, 64'h94630650b0d66e11, 64'h518c2ca6d7afb551, 64'h1660003e7b},{64'h6000000008040000, 64'hb13886e000005018, 64'h1036185934c859, 64'h3533c903f27000, 64'hf2a2663624c99318, 64'h18b660555a},{64'hc04018220000, 64'h6b06800000000014, 64'h9361c5c4c9879, 64'ha34bf65f554f41e8, 64'h119031f5a580c785, 64'hd07206258},{64'h806180050000, 64'h18800000000010, 64'h7c896b16fc54d600, 64'h5bc368698fce349d, 64'h15019446415107a5, 64'hcc00034f8},{64'h2000000146, 64'h24f6d40000000010, 64'h876b60505c5c9899, 64'hba1c76a06e00032b, 64'h9d8339a7346810a5, 64'hcf8dd3e56},{64'h2000000140, 64'h1c9a066000000010, 64'hc38f46185c456369, 64'he4aac112ab0460b, 64'h61981183f9800fff, 64'h19f0006d14},{64'h400000014000000, 64'h3159d24278003000, 64'h3b1788584c2cad41, 64'h9a1cf54ca999a277, 64'h189e164dc9358b9, 64'h70e0542e0},{64'h1000000106, 64'h1558d260b8000014, 64'h41b02e124c39e269, 64'hf035603800000405, 64'h8f8000708dfd835, 64'h7919562fe},{64'h4100050000, 64'h3116051210003000, 64'h7c492e264c2c8e79, 64'hab9e4dacca4fabe6, 64'h69adb6b1e0d6c075, 64'h83cf36b6d},{64'h8051902, 64'h3136800000000000, 64'h3cb6be24e4a96f61, 64'h13277c4dad53ceb5, 64'h4d14a154526a0d3b, 64'h130da0340c},{64'h1000000021800, 64'h1ca4840000000000, 64'hdad15cdf0c349861, 64'h62fad98c7239d0, 64'h11018e93e13a4d38, 64'hda36c41a8},{64'h104000c000000, 64'h309ba82000001000, 64'h978db3d6cc221899, 64'h6b4f35647d15a1da, 64'h6c0000056d9ca76a, 64'h106cee369d},{64'h400c00000010140, 64'h3140000000002000, 64'h5311be2d04ccb559, 64'he01f537d026aa28f, 64'h69ad6604336d4db0, 64'h13d7786b8d},{64'h4018200000, 64'h302bb4750800500c, 64'h540a5e233c3cd049, 64'hc7b47aab019964d0, 64'h450219740865db5e, 64'ha4d434c15},{64'h4000000000050040, 64'h160242000003010, 64'h554dabd9475c8b00, 64'h54578ae8d2668a85, 64'hceaa80035269caa9, 64'hd165b2a15},{64'h8030000, 64'hf014800000000000, 64'h3fd78e253c323073, 64'h4557ecfecfe41f, 64'hfdb0d4ae6c12b8, 64'h12b9b161a0},{64'h6, 64'h2ed5000000004100, 64'h38697e1c884d81a9, 64'h734081cff0f03f7, 64'h7cff9a43403f4d22, 64'h76d59bfe6},{64'h6000000008010000, 64'h1938800000000000, 64'h3e106e1f5c397255, 64'h201b1070cf84ae, 64'h92d89b0630c592b0, 64'h1839b15715},{64'h80000104, 64'h317acc0000000000, 64'h8af6861cfc25ac41, 64'h39c9e381268e0609, 64'h2d0580041ac59625, 64'h1063231c08},{64'h300000000020000, 64'hc5800000001010, 64'h97e1c8c4d5595, 64'h484be4ed375484e4, 64'hc8de66f0000009d9, 64'h12853b4b79},{64'h400000004000000, 64'hac00000000002000, 64'h158e2099b4985c, 64'h6d9aa878938270, 64'h492e672e30aa98b0, 64'h164cf15a6b},{64'h10030140, 64'h156a826000002000, 64'h56d44e1d00bc9859, 64'h3e553b216aec949b, 64'hf9b400027c521891, 64'h1667684c04},{64'h200000000030100, 64'hc4814180000000, 64'h99977e1cb8cc9500, 64'h502a000193f1f56d, 64'he079db86cededb39, 64'h7aa676406},{64'h1000004000080, 64'h1b28a6e810005300, 64'h534aa81c583cb859, 64'h3a409c5d82b171e9, 64'h8d8314b359c18a69, 64'h1b3eb8be65},{64'h100c000000, 64'h159894000000000, 64'hadcb8e20dbb28f00, 64'h1343769cf993e576, 64'he10921140b6a0cc6, 64'h9f800578a},{64'h865010200000, 64'h308aaeeab0000000, 64'hc14f9e1a5644b8a1, 64'ha0be3c1b0100065e, 64'h150b000377e6b005, 64'h138a8561ea},{64'h200000000000000, 64'h16a0000000000190, 64'h80cca6104c5ae149, 64'h5e29ac5d30000296, 64'h848c40049c859372, 64'h187f40c999},{64'h4000000, 64'hc609800000000010, 64'hd8948ae56c41c27d, 64'h5d40b57d66800578, 64'he15d26332c98d5e1, 64'hcb36329b4},{64'h803000000100, 64'h26f6a6ee40005080, 64'h3c1065964c519889, 64'h49e9347935a26f, 64'hcaf5b7093f5c0c, 64'h15e40f8000},{64'h40000000c000000, 64'h4400000000000014, 64'h129e2970bef86d, 64'he06b76a189996404, 64'h80a862b648981928, 64'hfa5b71e59},{64'h860014040000, 64'hb0f5867400000000, 64'h9b09ae1c5844986d, 64'hed625c4e6feb6332, 64'h6ccd00042b8a6748, 64'h80a6e3349},{64'h410001000000000, 64'h1000ea000005000, 64'hd6575a511c2acc00, 64'hb96b2000ac94d550, 64'ha4f9db49d3561025, 64'ha45491dca},{64'h500003010000000, 64'h31792eca08001000, 64'h1448aa5c3cb889, 64'hb53299aed2264000, 64'heca6f5a6b8aedadd, 64'h776656b8a},{64'h18004000000040, 64'hf5800000000000, 64'h654a6ba341548900, 64'h440865d022671c1, 64'ha5ae778b6a6dd31e, 64'hd18003789},{64'h20000040000, 64'hf110c8340cc00008, 64'h7d4bae1e8c389855, 64'h5787d4d1e5b574, 64'h9cd49f632f812fb0, 64'hfb25c2a36},{64'h1002180050800, 64'hb106800000000000, 64'h9ae2f34317895, 64'ha9cae44071ebcbf6, 64'hc06e800289c14aad, 64'hab705368e},{64'h10000200c0, 64'h30f4d85208004280, 64'hc94a2e184c2c9899, 64'hff348938fde4d1ff, 64'h108b2b3637fd2bd, 64'h6eda9e560},{64'h300001018442800, 64'h1af1825118000000, 64'h13ae186c5c9851, 64'h5740168382655e2a, 64'h58ffd9c33655c7ed, 64'haa19c2a8c},{64'h200001180042800, 64'h62bb000000000018, 64'hb2882a9c4c248d79, 64'h7c1a56ccd5539c0, 64'h30d8d4741aadd8c7, 64'h12c4e11db8},{64'h14040980200c0, 64'h161244000000000, 64'h4ed77e1cb94db800, 64'hdb57acc7053b49f, 64'h695915a1e5db0f86, 64'haa8006475},{64'h40000000102000c0, 64'h150dc2000000000, 64'h510b4366cc3c9800, 64'h6e6d74eea20004e5, 64'hc327000288554aaa, 64'h791552939},{64'h6000000004000140, 64'h4000000002010, 64'h3fd1661e9851d700, 64'h976314f8718df62f, 64'h4e8490832e3f9c19, 64'h155d49341b},{64'h1000020000, 64'h31174c2000004014, 64'h440dab1f4b813881, 64'ha06ce68164d002a0, 64'h80a80e06403b09f5, 64'h1b655cc1b6},{64'h18001100040000, 64'he6e0482000000000, 64'h37576e2ccc55f88a, 64'h7ba9ac187d54b290, 64'h25905b8d56aa5b3f, 64'h1548de5945},{64'h500040000060000, 64'h9baed310004000, 64'he7e2550a91800, 64'h3503e5555b0588, 64'hc5305b12c7c1b618, 64'ha6cfb2e66},{64'h118800000000100, 64'h7009000000005000, 64'h9b1686133c2ead51, 64'h4e66dcff2a74d1, 64'h4d095f4c29934000, 64'ha1ea83488},{64'h6400002000000000, 64'hf09a800000000004, 64'hcf4ba626ac5c9893, 64'hd42dc359e8004c0, 64'h172ddfa3f400198f, 64'h12f9fa4e3a},{64'h410000000000000, 64'h2e0000000000100c, 64'hd4bac804493a1, 64'h5788215d15d000, 64'hb586e70c10ab5568, 64'ha753942fa},{64'h400010000000, 64'h4600000000000008, 64'h464f5c25403893aa, 64'h5b40fd6d270001e4, 64'hc95f8002719387eb, 64'h8d2bf59d3},{64'hc00014000100, 64'h10c4c47318000000, 64'h6d947e2cb0c162b9, 64'hf058982d27d951f1, 64'hfd162296b78b1059, 64'h1042bf410a},{64'h4400001000000000, 64'h46b4a90000000000, 64'h6557ae2049b08f6c, 64'ha73527c8dc00036c, 64'h8705e5c3346a592d, 64'h1369f336f3},{64'h200000000000000, 64'h40e1000000000004, 64'ha996bd133c3e3243, 64'h54cafcaeada494, 64'ha8cd5392b24e55f8, 64'ha1a4b203a},{64'h400000000c00010a, 64'hf1385e49b0000004, 64'haaae401a47d098aa, 64'h63739ac00000271, 64'h6726000648c19b43, 64'h130a4c29d5},{64'h400005080060000, 64'h30c4c5e000002000, 64'h82e265c38d881, 64'hb6b469a98966a40c, 64'h1db46076b93f5305, 64'h132cf11fc8},{64'h1190400000, 64'h6a00000000005300, 64'h3c8bb3432c3d2a99, 64'hbdaa16db01800424, 64'h7134cf31e4858dbd, 64'h133cf5bec9},{64'h5000040080, 64'ha0816000001180, 64'h9a0fa62ee6d8b800, 64'h4027e0018bec8353, 64'ha02694d252cf9d, 64'hfb6bda960},{64'hc000001180000000, 64'h22f5000000004114, 64'h938dbbaa5c489861, 64'h14ca253d2894f369, 64'hf2850e04a253c6ed, 64'h9fd0cd71a},{64'h218400000000000, 64'hb800000000010, 64'h6acc6e26fac9d400, 64'h581da4dc9b9ab1da, 64'h8d9372bc255618c1, 64'ha680061fc},{64'h200003000010000, 64'h317ad26000004000, 64'h16961e88c09859, 64'hd4bc4bccde6425e, 64'h34ce4006c8978abe, 64'h18c6b82a98},{64'h10c0000020000, 64'h3169c9e000005000, 64'h9b9158409c38b8a9, 64'h5a33cb0cadeb2588, 64'h155999e4c765acf2, 64'h1b1ecbd66b},{64'h10080, 64'h5800000000000000, 64'h98178e2d35c1b255, 64'hba2aa64d59f266d9, 64'he8ad66c57464d359, 64'ha29a74bea},{64'h1001000053080, 64'h7137b96814820000, 64'hc2175620a6d4d88a, 64'h6b4ddb3cd4713a89, 64'h51849544c1ad8aae, 64'h12f8006125},{64'h400c000044, 64'hd5800000005000, 64'h572abb228c4df800, 64'hf707c3cd037f1ff, 64'hd484eab1ea00074f, 64'h15bced61e3},{64'hc10000000c000104, 64'h30e5d06000000014, 64'h403154c49c34b8a9, 64'h341aaca6abb6b3, 64'hbaa8eab229ac5588, 64'ha6aa95533},{64'h1000100000000, 64'h107800000000000, 64'hd88d4ce880d49800, 64'hcad840010c2c241e, 64'hd47a8005776c555e, 64'hdf8006c63},{64'h6200004014e60000, 64'h70c5d64abbc40004, 64'h4dd636107c5098a1, 64'h1340965f025f7206, 64'hd6d8f131e0ebd027, 64'h162df81f75},{64'h4000010000, 64'h1200000000003008, 64'hcb4fbe2cec45b8a9, 64'hfa34ec08dbf0d65c, 64'h1909e60352c08fb5, 64'h13ae614ddc},{64'h1000018400146, 64'h2d37c41510000000, 64'hcf6e9612d0ac98b9, 64'h4afc375e0fa3f7, 64'hbc7d9ef60b7eb8b0, 64'h15e3231f67},{64'h1006008600140, 64'hd5800000000000, 64'h9389861556510100, 64'hadc1157ed4255349, 64'h58da1f63ff7d8ffe, 64'h198a563689},{64'h8000000, 64'hf682e000001190, 64'h9aad546209800, 64'h241fbacd05b13566, 64'h8800df56400192b, 64'h79d1ae2d4},{64'h800004000106, 64'h140800000005000, 64'h8b2c6ae3584dd600, 64'haf4174f0d416b1c1, 64'hecdbd3c4596bcd49, 64'h70d3a3e64},{64'h40140, 64'h117854000003000, 64'h7ed55e2141353300, 64'h8c27295c9ddb8a77, 64'h60fe08c56c7f09c8, 64'h1376585b89},{64'h400400000000080, 64'h116c03208000000, 64'h3a499ad977a9c300, 64'had55ab28ad5952bb, 64'h796b627366074a, 64'hcc0ea0000},{64'h240144000c0, 64'h128800000000000, 64'hae936e1157de0900, 64'hfd27dc96db9a46d1, 64'he8792c74c39b2cbc, 64'haeac82b64},{64'h1000014030000, 64'h400000000000000, 64'hc14dba54b452a18b, 64'h366cf565354e0204, 64'hd103f746413786f3, 64'ha40f31c2d},{64'h18020000, 64'hf0d5aaa148004014, 64'h51d3461e4858988d, 64'h6960db210a55b2b8, 64'h45092073fe81d0b6, 64'h6f6b72938},{64'h3000000100, 64'hf6c40000002000, 64'h9455bd96e64d2100, 64'h9359caa9662e0351, 64'ha9541aa4d364ca05, 64'ha06ab59e6},{64'h11000, 64'h30d5a6717dc44000, 64'h690c2628492898a9, 64'hb536c000a7e51a17, 64'h158c20540a80d021, 64'h1544ee62c8},{64'h10000000c0, 64'h8404800000000000, 64'h83cb7e2379360e62, 64'h427cc810695a647, 64'hbcacb1f2b07bcac6, 64'h10815929a7},{64'h2000000046, 64'haaf5d00000000000, 64'h992e5266dc5e2864, 64'hc041bb10cf2c0597, 64'h89ad362566c99b26, 64'h162b126fcd},{64'h418005018400000, 64'h30d5b87410000000, 64'h53cf4e1130c49553, 64'hc06b767aa78fe57e, 64'hb55feb3cc0001ade, 64'h137e615803},{64'ha1000000080000c0, 64'h317a000000000010, 64'h6e555e12e0588a89, 64'h64f9ad64ac8375, 64'h2336660612b1d638, 64'h15c2bc57f8},{64'h1000000020000, 64'h30e0000000000000, 64'h39cf4c2a8a4da1b9, 64'hb11ce0016870f554, 64'hb984c00335d6955b, 64'h7435a2023},{64'h10000140, 64'h70f4d4000000600c, 64'haed79214b0c2c289, 64'h4c57fc3f8200054d, 64'hf49e800556c1d54a, 64'h125f077034},{64'h400005000000040, 64'hc58ae000000000, 64'hc809a3dd00449800, 64'hb6640814a6a0429b, 64'h126605334c7d835, 64'hda94e29a0},{64'h200080, 64'ha200000000003000, 64'h6a4dace4fbd14943, 64'ha94216fef9943431, 64'h14295e49a578f89, 64'h10cda93e80},{64'h101400000000004, 64'hb000000000003010, 64'hc4edabe29bd20a63, 64'h9863065cb8b172cd, 64'h80825984b9c198c1, 64'hfc5393ed5},{64'h10000000000c0, 64'h7027800000000004, 64'h988b4e1b38c2b2a2, 64'h514c46e8d4f1765d, 64'h8c840512973ec6f8, 64'h1319a84c3c},{64'h100000000000080, 64'h4116bc2000004000, 64'h6b0c86269c5e485d, 64'h6b3585ac79000579, 64'h9c7de566e879cae9, 64'h127cf16e87},{64'h100000008050100, 64'h66f5b94d00000000, 64'hc4d44e244bc0b889, 64'h31663c4c9bf05357, 64'hc4da4e0200034981, 64'h19300d4ad4},{64'h1014000104, 64'h22f4de6000000000, 64'hace8ae1cd0409859, 64'h3a4bd9b95e26e25f, 64'hf00000027851d92d, 64'h15ea4f2daa},{64'h4000000, 64'hc000000000000000, 64'hd9934d68b43a2253, 64'hbc353d65d8359326, 64'ha2a5828a000fe2, 64'h6ce0},{64'h201420010e00000, 64'h30abd6700b406000, 64'h93cc33a25c5898a1, 64'ha9327556d4a4f350, 64'ha96f4005757f2ab9, 64'ha2e4f4b13},{64'h400400000000000, 64'hb1000000002000, 64'h3d954de36a409800, 64'h1ec3d5654f5276, 64'h88aa5a233156c000, 64'h755a13426},{64'h1000008050000, 64'h5b5980000000000c, 64'h81892a9f60c89759, 64'h7d371384d05591c2, 64'h243e8001eb845088, 64'h1644e11fd5},{64'h4080000000, 64'h116000000002180, 64'hfbc269b556000, 64'hdeec83d9083631ba, 64'h798d8006c8c6d58c, 64'h81f3abec3},{64'h401c00000050004, 64'h30f62ec000000018, 64'hb274506a6c38d299, 64'hf11be849614e12b9, 64'h407ad08363aec709, 64'h6c7b},{64'hc00004000000, 64'hc400000000000000, 64'hcf4d96271c42555b, 64'h359d8118d303604, 64'h102b285c9ca9547, 64'h18da524a40},{64'h8050102600c0, 64'hb0a4d628a0000000, 64'h928c982c4c348fb9, 64'h1c6056db86d58631, 64'h2caa00040b870fd6, 64'h10aa234469},{64'h400000000011800, 64'h14bb800000002000, 64'h3f9560104c3c9149, 64'h144247c59055a9fe, 64'h38f7ec549c52ca6a, 64'h10867f1dc5},{64'h2001060000020000, 64'hb0d0800000000014, 64'h38d29c60f5dd564b, 64'hb157e555606b1562, 64'h16ad0003eddfb936, 64'h1600e449fb},{64'h10000000c040000, 64'h9b800000000000, 64'hc9e2b1b224200, 64'h5817c905daf35e, 64'hb930e23424970ff8, 64'h8066d4229},{64'h1404000011000, 64'hf00000000000000c, 64'h7c497ad50754966c, 64'hc7c346b164e6baba, 64'ha16aa523e7ae8d7e, 64'hd62523773},{64'h4298020000, 64'hc6d4ac0000000080, 64'h935346257c58d863, 64'h39a7393955db1362, 64'h6182996362660465, 64'h74502e0e6},{64'h10220000, 64'h0, 64'h8153be16d7d5d653, 64'h2955baaf2672029a, 64'h84dba61640814cbb, 64'h18b20636e9},{64'h3000000000, 64'h9bb562b01e0000, 64'h371146150655c100, 64'hfd352a986e2a63e6, 64'h1bab191e4510db4, 64'hf93756320},{64'h430003000000000, 64'h18d55677a0640014, 64'hc61640a2ec01f849, 64'h102aa00134a0f4d2, 64'h59ba4f3abd80d446, 64'hab0001c35},{64'h1065088000000, 64'h171000000000000, 64'h64d57c5125d0b600, 64'h98e31700e00002c3, 64'hb0dcaac40f5d734d, 64'hca0e14c6a},{64'h4180060000101c0, 64'ha8d5a84000005100, 64'h4dd732186c013899, 64'h6b6f6000dd5ac4a3, 64'hd5723a116b0c9d, 64'h155e63ed00},{64'h400000008600000, 64'h0, 64'h4ed1be24ac55e100, 64'h1e2bb5ae9e000760, 64'h387753f63c4fc9e3, 64'h1072231e78},{64'h2001003000050000, 64'h30f6c5c000002000, 64'hd950bd1055d89849, 64'h3c4d6dd506d3b578, 64'hb363743df98098d, 64'h98f6664d4},{64'h419400000060000, 64'h121b000000000000, 64'h93536e24f646a2b9, 64'h6c49e000cf66eca2, 64'h8db156fd674e8a2a, 64'he126e34e5},{64'h4000000000000100, 64'h8700000000000004, 64'hacd2be16fc46c942, 64'h352ab559ac929f, 64'h53641ad28baccd68, 64'hd600057b6},{64'h1000000000000, 64'h19000000002000, 64'ha9cd44193ad1f700, 64'h232b6aad552a749f, 64'h6cd082361351d558, 64'hac710620d},{64'h301000000050080, 64'h3116deac00000000, 64'h3f90a4d25549e159, 64'h6827a5a187c001ed, 64'h6cd14ee6b5b1c9e9, 64'h8019b3436},{64'h428000000000044, 64'h26b4800000000000, 64'h56b76a1e5c409289, 64'hb657cca4cf2be1c3, 64'h9eebcd7c3c508d, 64'h8231736a0},{64'h8030000, 64'h2200000000000004, 64'h84934e10fc49d555, 64'h6c93847b53b1c0, 64'hbd095f321056cad8, 64'h1b78006c9d},{64'hc0, 64'h80b4000000000000, 64'h840fac27615da175, 64'hfa6e8001b1b745a1, 64'h590900040ac15949, 64'h1b236360ec},{64'h400c0, 64'hc55901c000000004, 64'h53d44a2f1629f882, 64'h631f6561834fb67f, 64'h74ce800612d8d92b, 64'h293246076},{64'h6001404100000000, 64'h30c5c5e000000004, 64'h848974245acee041, 64'h1cbde984f7a6129a, 64'h8ef78001f77cc28e, 64'h1ba9e842b8},{64'h6010a3000000080, 64'h315986c000000000, 64'h3c92652ef020b849, 64'hd722001c22ad1ff, 64'h12b4f23cfdd3414, 64'h1592ae1e60},{64'h1000000000142, 64'h309aa02000000008, 64'hac776aa24c509891, 64'h5164ec4927951627, 64'h3ca800001b56b931, 64'hd82505819},{64'h400000030080, 64'h81000000000000, 64'h7f11656139516900, 64'h44b0869135fc35f, 64'h2802000425d9d2c0, 64'hf930a4ddc},{64'h7000060000508c0, 64'h31162d2000000110, 64'h939535e0793c989a, 64'hea2749b9ace1adab, 64'h3d2c6701d44ecfe4, 64'hd6d60ecf9},{64'h460000000080, 64'hb800000000010, 64'h6a135b5f2c389100, 64'hc202844da211363, 64'hd07b0f5331c1e80a, 64'h1908f61d56},{64'h100000000040004, 64'h2481000000000000, 64'hc8338d577a25ac81, 64'h24bcc0c7ae60653, 64'hdbdf34c2c0981b, 64'hfa1450fc0},{64'h118004100000000, 64'h3117ce0000000000, 64'hc6d59390d0093851, 64'h5ec084098d90441e, 64'h7f7759bc1cc3ed, 64'h1350dd0e60},{64'h2001000000000080, 64'h6af5204000000014, 64'h6c56901c5c50979a, 64'h6c6d87d0fa0004d3, 64'h5aca198637660cbb, 64'hd936c1bd5},{64'h400000030000, 64'h149a2ec00000100, 64'h98d14c9b07800000, 64'h1c636d9ce06634a4, 64'h598e156373001bdb, 64'hca509ca65},{64'h50880, 64'h157ab56000006010, 64'h80d236213c30d1b1, 64'h4b42a7d581f7bb59, 64'h95070002df92d0aa, 64'h18de4b4a58},{64'h2000800000000000, 64'hc6c0800000000010, 64'h658f4c61393c985d, 64'hf58add49e5b86ea, 64'h3a2d00f43ddd1628, 64'hdb85a4978},{64'h408000008000000, 64'h116b12000003000, 64'h38137d917ac09200, 64'h4e279401bac00276, 64'h6d62e6c9ca538801, 64'h1b366f4e09},{64'h10000000c000000, 64'h3117800000004100, 64'had90bcd2b506d871, 64'h3854f09e2ca596, 64'h90b1e134287fd318, 64'h7266eca19},{64'h10080, 64'h149800000000000, 64'h948b862b7b35ee00, 64'h1a00000164d5b567, 64'h51881186b6c68d6f, 64'ha41946346},{64'h2400000000000000, 64'h70b4b02370000014, 64'hc5cf546a815c9869, 64'h115579b09eb18566, 64'h432965640e0018c2, 64'h15a26e1d1c},{64'h8600000, 64'h8b504000000004, 64'hc5d176217acda900, 64'h927b5a38480057c, 64'h34792724c0af55eb, 64'h8055f5915},{64'h50000301c001000, 64'hf148c1f610004304, 64'h95e02cc35d805, 64'hcc40b40994ebe9c2, 64'h5d30cdd1ba658db6, 64'h10354ea096},{64'h40000018005098e, 64'h7160800000002000, 64'h6a6b7e1a674cd889, 64'h8e04935534e19b9, 64'hf98cf364ec000add, 64'h109d5e2bc4},{64'h100c00008000100, 64'h0, 64'h3ece9e12b5365800, 64'hac60fab186800631, 64'h1096e1655b84ac2, 64'h1b254e6480},{64'h400c00000010000, 64'h1f70800000000014, 64'hc4d0489540449369, 64'h556c947deab3fc, 64'h4d565f40a57cd920, 64'hf81f44c78},{64'h803000000000, 64'h159200000000000, 64'h5650bcd2f6aec100, 64'h3f67e000f7f1e63c, 64'h9cb61e76eb53cf47, 64'h7995a2d87},{64'h104500c000040, 64'h18d5810000000000, 64'h93d77a6a5b44b251, 64'h772dc187e80001b, 64'hf98380027fe1f8f7, 64'h1670f55783},{64'h4000000, 64'h2b800000004000, 64'h3e0c9c6895a15800, 64'hfe64f000a8e581fe, 64'he47ca714e2945b38, 64'h15edfd1d03},{64'h4004000006, 64'h90542280000000, 64'h86ad7b9776455600, 64'h64b13a95e2c23f9, 64'hd5e30760e3d4a2f, 64'h1618f657ab},{64'h2000040000, 64'h1531000000001000, 64'h97e1155b62ea3, 64'h9a356668d4cf5358, 64'hd9386a8368aa0755, 64'h9e5ad41a3},{64'h60000400c000140, 64'h5f38a6c000000000, 64'h71ce9040ac2ea269, 64'h452036d508db554f, 64'hacd0e674ce00011d, 64'he42674c26},{64'h2000003008000000, 64'h1005000000000010, 64'h6a535d5a970a38b9, 64'hde2bd4ed5935a368, 64'hd2da2cd59a0003f4, 64'h9e37b3377},{64'h30080, 64'h89862000000000, 64'hdb09ae1b4732f600, 64'h986f298882779637, 64'hb5cda6d736b1d085, 64'h1640005789},{64'h400000000000, 64'h1d10dc0000000010, 64'h874b9b5ea4489561, 64'hb66d9811b78006f2, 64'he0da9a13310e10b1, 64'h1bd3706df0},{64'h5104040000, 64'h70f5a6800000000c, 64'hc6c613c5888b9, 64'h1cef9685ba5a1704, 64'hd8000006dadad02f, 64'h18e7834a77},{64'h4000050040000c0, 64'h2a20000000000000, 64'h6d4e7e02bc58a999, 64'h4bc2b65d629b044d, 64'h88cee8750e001b1e, 64'h1311b636e9},{64'h8040000, 64'h1d41000000000014, 64'h8557aa5530a08b69, 64'haf58bab930e156eb, 64'h85579fb000000802, 64'h29d3},{64'h3000000080, 64'h2200000000004284, 64'hc5d56de0bc4c9861, 64'hca2013f5553232c7, 64'h8c7f0f359400072e, 64'h1576b2ce1c},{64'h800000000040, 64'h4000, 64'h56cbbd5d48cdac00, 64'h4863462c02a6b597, 64'h193626142962d325, 64'hd840000a0},{64'h218004000000000, 64'h1737c80000000014, 64'h6e956b2f10a898a1, 64'h1ae309b8dd1a849a, 64'h7d29d1acee9d8027, 64'haf94d6155},{64'h400000000000000, 64'h9c19000000002000, 64'hc114add095cc987d, 64'h5e42081593b5e64a, 64'h127f21642c89913, 64'h1376104250},{64'h402000000000, 64'h2158800000004180, 64'hcb56bd1339348e79, 64'hdd1bacbd9793e27c, 64'haff2820965d394, 64'h190f2ae0a0},{64'h404014620000, 64'h16a81f10c820000, 64'hc617561a4c4c9400, 64'h83607b3281483646, 64'h5d918ba1bbce1814, 64'h3a0ba49ec},{64'h1000000000000, 64'hc4d4d62000005004, 64'hcbd80ac20987a, 64'hf34b43cd561c04dc, 64'hd4d92700e76c93b4, 64'h1355f52bd7},{64'h600c01008040000, 64'hb138d04000005000, 64'h6596935857a48ba9, 64'h56559558fa537380, 64'he0ca5385c356992d, 64'hd9559be84},{64'h500002000000100, 64'h7015000000000000, 64'h53d6be1756c4b379, 64'h5864b0016493b4c7, 64'h38ab56359058d0a5, 64'h18fab22b25},{64'h418000008000040, 64'hf080800000000000, 64'h168dabe2b5393405, 64'he467f03c2d80063d, 64'h10756cd523902d8, 64'had4105a40},{64'h510004000000000, 64'h1317800000000004, 64'h538a762e5c40b499, 64'h7800000a72074a2, 64'hd02d6ce9f282007f, 64'hba0001fd5},{64'h100004000000080, 64'h16e0800000000000, 64'haf0fae016c509741, 64'h72a04e8000001ff, 64'h447cec34e34f0a77, 64'hb91512745},{64'h40000040000, 64'h3bb43110000004, 64'h8561f3c264b00, 64'h9f55064c9e5a96b2, 64'he8da1c71edc1f541, 64'hdd35c5876},{64'h510c00000060040, 64'hf101c86000000010, 64'hc909b61115b2a06c, 64'hb527c6adadf1f423, 64'h79884f6d51ad533a, 64'h1928003295},{64'h400000050000, 64'h2300800000004180, 64'h17aa1721027879, 64'h96d0c249edb5b56, 64'ha1659ad4cfacdb43, 64'h15a5c8d96d},{64'h405000040184, 64'h5938800000000000, 64'h6d2db620b905f851, 64'hc760e00184f0657d, 64'h8d5a30759bad15ee, 64'h15eab46f79},{64'hc00000020100, 64'hf000000000000000, 64'haf8dac9897c50102, 64'h4536c651bcd5a1c3, 64'h5536cff7373fcac9, 64'h1649951f46},{64'h10000, 64'h6b20000000002180, 64'h38c99ad17c354f84, 64'h6b6dadad0b60d422, 64'h90818e36da000db7, 64'h1bd61ea063},{64'h30102, 64'hf0bb800000002000, 64'h85aa6b2d5c3a3274, 64'h1c25e000d0d2f1f7, 64'h553101f36e6c5b6e, 64'h1c1c1f3468},{64'hc00000040000, 64'h70d4d64c10005008, 64'h3a0e5040fc2cb889, 64'h33d035155cd43f6, 64'h19231050f40d929, 64'hf85b6cc50},{64'h400403000000000, 64'h3159800000002014, 64'hc68fbc58d802d891, 64'h60000018d30642b, 64'h98f3f26205b2957f, 64'h157eab1e7c},{64'h200001000000000, 64'h17a000000004000, 64'h350bae1716bd3800, 64'h5b1a829591d3c4d6, 64'h247f6c96f2295655, 64'h1286c44c6b},{64'h8053000, 64'hb137de400000400c, 64'hb4b6350d94071, 64'hb7bd2c767800, 64'h9278f61ec7bd3b1, 64'hfece100d4},{64'h2010000000, 64'he6800000000004, 64'hc1537e2295c18300, 64'h211d566c00000375, 64'hdc2ae336ab9387, 64'h19319c2bf0},{64'h803010200000, 64'h70f6c44000005000, 64'hd748b81c49a49861, 64'h3358433f35d65a, 64'h182a4c6439cd914, 64'hd6e854960},{64'h1020000020000, 64'hb17a800000000000, 64'h3fd6661edc25b8a2, 64'h51fc3a997c0022c, 64'hb88e36e4c3ca3082, 64'h1976101bcd},{64'h6000800014000000, 64'hb0d5800000004004, 64'h65498c253bb0b8b2, 64'h6d1bde0d371cd647, 64'heafaa680e99b4d92, 64'h9e6504efc},{64'h300404000000140, 64'hf100b04000000008, 64'he0f6c68904cb8ad, 64'h716e0c90ab3246d9, 64'h68e1f713654e0cc7, 64'h3ebc},{64'h101000188000000, 64'h31413c2000005000, 64'hc2135d645c34b1b9, 64'h5aaad001d7b28650, 64'h609c68a071658e15, 64'h1b84004966},{64'h10620000, 64'hb000000000000004, 64'h7ccb7e2b7b3498a2, 64'hff49756b64f59554, 64'hc90984b2c7d710a1, 64'h1ae04b2b37},{64'h8000000041000, 64'hb0d4800000003000, 64'h6f975e1157b23005, 64'h41fa85962c5bb7e, 64'hcd6945bb2c0010b2, 64'h854f1fc3},{64'h4000080, 64'h9100000000000c, 64'hdad775a119c96a00, 64'h484e581d0466b29d, 64'hb0a89734d89849e1, 64'h9e2092e9d},{64'h0, 64'h40bbb04000000008, 64'hab499e2af741016c, 64'h526b6949568006d4, 64'h81ae18c000000da2, 64'hd836b2a36},{64'h6000000010a00000, 64'h3138de89b0000004, 64'h7d904082bc324069, 64'h317c6b0d1f6434, 64'h2f091f3640db1b58, 64'h1089fd3757},{64'h443000040000, 64'hb17a800000000000, 64'hafd46d9f0c212c03, 64'h286060018c7686d0, 64'hc8822bf2bf6db5af, 64'h192eb42083},{64'h300002004040000, 64'h7150d82000000000, 64'h6611962edc296c12, 64'hb46d1b1daf50257c, 64'h7d65d4035bc1d66e, 64'hccb5f36ed},{64'h40601c050106, 64'hf0b4a2f1081e0000, 64'h9b73b0945c3498a9, 64'hf41bbc0ccbcfa27d, 64'h10ca8845696546ec, 64'h7fb041fec},{64'h400800004051800, 64'h70c03c0000000000, 64'hdb099ad1150ab869, 64'h715939c441d5a9e6, 64'h5d5011ff405b6a, 64'h7a25732b0},{64'h10450000, 64'hc600000000001000, 64'h114cec44348f85, 64'h511e7db75661a6d4, 64'hac81db73e6000cc1, 64'h1095b22a0d},{64'h400002000000000, 64'hb0bb000000003004, 64'ha991561b000538ab, 64'hfc64a7a0ad0e32b4, 64'h9cfa5033ce0010bd, 64'h10fde936da},{64'h800000c0, 64'h936a482000004100, 64'h270bbe1b5c0a389b, 64'h25d5227191b183d1, 64'h6888b23222aac81f, 64'h18fe16efcd},{64'h110004000000000, 64'h1d79800000000000, 64'hdbcf9614bc36b461, 64'h8588820f836f3e0, 64'h21936ccbe0000726, 64'h19455c2928},{64'h1100000c000000, 64'hb17a800000000000, 64'hc11475a2b9a54104, 64'he96f5400f78001c2, 64'h3164e6c9f356c818, 64'h9e18c6566},{64'h500806000000000, 64'hf0b4828000000010, 64'hf46211c4ec155, 64'h3960c57d362582ba, 64'h9961c004efdad83d, 64'h13737857bc},{64'hc04014200000, 64'h8000000000000008, 64'h168cd2fc52a85c, 64'h655166f3513c2c6, 64'hb13600037158d547, 64'h19726a3399},{64'h4008600000, 64'h3000000000000004, 64'h79cfad96962220a1, 64'hf0511a0af3800230, 64'h413926040e9c933c, 64'h8030b4eb8},{64'h800010000040, 64'h477a202000000000, 64'h9a0c6bd6e02498b4, 64'h5e613d78000001ff, 64'hf52d9a423900163b, 64'h1379cf590a},{64'h80, 64'h4738800000000000, 64'h65905a90c082f84b, 64'hc76349512a000707, 64'h7d0715f00000136d, 64'h10914e4245},{64'h300002010000000, 64'hf149800000001000, 64'hb4b50c502588d, 64'h36d39592597000, 64'ha41cd98612395b8c, 64'h1b8ecc594a},{64'h6000002000000040, 64'h2600000000000010, 64'hc1ca5a42ec36a079, 64'h5b0402700f89c651, 64'heafa35c040001457, 64'h109b081c99},{64'h4300000000500c0, 64'h2559a6e000000000, 64'h3f48609b10d09871, 64'he61cc00097d975a5, 64'ha40fe62be93e5870, 64'hdfb291acc},{64'h4040000, 64'h3128800000000000, 64'h982eef122a051, 64'h4142d4f06a607000, 64'hb504b1c4a0505281, 64'h104acd59aa},{64'h300400000000100, 64'h117c1c298000000, 64'h7e08ab12b5349800, 64'hd653c1a8d029e635, 64'h58baca64d91a86a8, 64'hfc8004133},{64'h100002010001940, 64'h6337d648b8000000, 64'hd8c1a6205c349859, 64'h6314bdb0da58c9a9, 64'hdd4e2424389ae7, 64'h190b640000},{64'h201000000000000, 64'hf6b8419800000c, 64'hab978a468c000000, 64'hf300000157270435, 64'h1094001ed7d1911, 64'hfa24b64bb},{64'h201005000600000, 64'h7015800000000000, 64'h154e1117d09781, 64'h97651b37639ba350, 64'h5c826c355d7bd90d, 64'hdfa1537e8},{64'h800000000100, 64'h400000000000100c, 64'h90897aeb6c222aa3, 64'hf06dc970f825c6bb, 64'hc000002813edb71, 64'hdccf520b9},{64'h240000200c000000, 64'h2559aee000000000, 64'h148e04fc053881, 64'had10995d94b17652, 64'hffb760635a8187fd, 64'hd6a066093},{64'h500804000030000, 64'hf000000000001000, 64'ha78d4be95b391104, 64'hb74e3a79b6da3434, 64'hfadf4203d68d95, 64'h7a5776b80},{64'h201400000040000, 64'h7179800000000000, 64'ha7e2350d9a349, 64'h8b2a36d0ab5b46ba, 64'h78db75e27162cd91, 64'h1672bc59cd},{64'h1000000000, 64'h117800000003008, 64'h804bb350954e1500, 64'hab634d6d00800096, 64'h94d280054fc8c826, 64'hf4eab42d6},{64'h408c00000000000, 64'h317a316000000000, 64'h908f90a2900678b1, 64'h7a2b4d9d041562b0, 64'hd025f7ea23de4ad3, 64'haca433e25},{64'hc00004000000, 64'h309bd02a00004100, 64'h1b8f9c61595aa859, 64'h6c4111b8803743e1, 64'hd5bab70593dc0763, 64'ha7d5d9d4d},{64'h500003004000000, 64'h3179bda000000010, 64'hd70bab2901055889, 64'he1207575cd0df734, 64'hb8a8d5da70e0d964, 64'h1ae8006d99},{64'h10030140, 64'hac8bac4000006104, 64'h11ae26e03cd8a1, 64'h734a588d93e2355b, 64'hdd62800592dccfb3, 64'h1b5e6eef17},{64'h118000000000100, 64'h117800000000008, 64'h58eb861ccc4c9500, 64'h764989d9818003ed, 64'h313666bf34001262, 64'h127b0465d9},{64'h1180040140, 64'h3000000000000008, 64'he209a62289c17271, 64'h1ad9a1b9b446e6d1, 64'hd137b2b4e5971085, 64'h1c48f46173},{64'h601c400000, 64'hf159ad2000005190, 64'hc78646c5c8869, 64'hcd60f9b6ca1d2376, 64'h22ca00037274d5a5, 64'hccdd1ebfb},{64'h401440000000000, 64'h3000000000003004, 64'hde8e662d4c558f8d, 64'hb44387c964b5942c, 64'h58cad5fb2bc97642, 64'he5dfd4258},{64'h8600000, 64'h6800000000000004, 64'h21d29e2f5c2d3684, 64'he3313972788772e, 64'h41b6a4f426001ae0, 64'h1666006559},{64'h400040000c000000, 64'h717ac02000000010, 64'h62546adc903098b4, 64'h690419b4c48001f6, 64'h83360006b957d33a, 64'h7f26c6d70},{64'hc00014000104, 64'h317a000000000000, 64'h6ff38e130622c179, 64'h564b85905a162b5, 64'h984f2101ad275082, 64'h4f1a66536},{64'h800000000100, 64'h18b4800000000004, 64'hdc138d5b483c9841, 64'h536e066082102139, 64'h4904f716396606ea, 64'h59b9},{64'h3008000100, 64'h3137800000001000, 64'haa915e2b0a489769, 64'h2e14d544a8aa66df, 64'h9ca8aa7375b286b6, 64'h6b6cc6c8a},{64'h100000000000140, 64'h70a0000000000010, 64'hab4bab66ca3ee989, 64'hbc55cdf1bdb683df, 64'hd192db636c6f0d91, 64'h1b25a33197},{64'h30000, 64'hc415800000000000, 64'hb1cf4c6959b60e95, 64'h9b336001916c54e1, 64'h6cd0b25374c95909, 64'h3766},{64'h4000000000000000, 64'h4600000000001000, 64'h7c115c9b07b98abd, 64'h5c2a0001b73271f6, 64'hfef3b263d0571839, 64'hddde842f6},{64'h4600100, 64'h1c0bd06000005000, 64'h3d8f945b0a86c24b, 64'haf1ffdba7b0af3cf, 64'h3d2c1301ec4c1030, 64'h80760652c},{64'h2010030040, 64'h3158bdb000000000, 64'h281475d4bc0d9849, 64'h396bd6dd38f5b653, 64'h54d235c40d000d6d, 64'h12a8a12ee9},{64'h800000040000, 64'h169b800000000000, 64'h6e93605b502a2341, 64'h9835a6fd2a5a9368, 64'h90b1800437d78d69, 64'hdd93c37e5},{64'h20000, 64'h128584f00000004, 64'hc4aef542a3300, 64'hde556274da4de140, 64'h85af708610275918, 64'h18f89e59d2},{64'h300000000040080, 64'h3158aec190005000, 64'h3990401a573c9349, 64'h626c40004e7686fd, 64'h90267624c898dbcb, 64'h1844e72b29},{64'h102000c0, 64'h12a1000000002000, 64'h40116c96f742a0b9, 64'h1cd56b5524b2eb, 64'h39692ce6eab49258, 64'hacebd1dab},{64'h4280020180, 64'h158380000003000, 64'h800b4b5947dd4100, 64'h509c200081d5e279, 64'hadbadf92967e4a0e, 64'h1b6e011c21},{64'h100510c0, 64'h309b800000006000, 64'h85d2502ae0b4cf59, 64'h170d57c54f783f35, 64'h388200e22e411149, 64'hfcc001e60},{64'h10a0080061000, 64'h22d5800000000000, 64'hab4c53ef3c427871, 64'hc9edadb1b6623c98, 64'h1b6aaf1c584afbe, 64'h1b5b6d6080},{64'h400000004400000, 64'h9981561000000c, 64'h568dbe1889000000, 64'h4ed932721f72b8, 64'h91606614e47d9390, 64'hae8007393},{64'h4000000000c0, 64'hd000000000002000, 64'h6f157e28bc39b0b5, 64'h37293121a4c659, 64'ha13853859d6549c0, 64'h1c4e5d4ba6},{64'h6000800000040000, 64'hc306d66000000014, 64'h4f142e24f0248aba, 64'h5b1d40012e503592, 64'h46ae8003a7848821, 64'h10ea004877},{64'h100000000030080, 64'h4161800000000000, 64'h93d1bb2b2809f842, 64'h9f400ab564f9a42d, 64'h35bdd4a59c52909a, 64'h6d6b},{64'h104, 64'h86f682e000000000, 64'hdb6b9ba120c498aa, 64'h553189d84385553d, 64'hbc7f18c4d8dbdb78, 64'h1280884eed},{64'h100004180000000, 64'h158a68c13820008, 64'hc68f5c2685349200, 64'h5fe36c1936c00636, 64'had3660e420000c5d, 64'h115b2e1fd8},{64'h518000000001100, 64'h1600000000000000, 64'h40899e257b39a141, 64'hee1dc0010b49dc03, 64'hbcd2c9ec888a5170, 64'hf80001bc8},{64'hc00000050080, 64'hb128800000004018, 64'h5457505c4c410b79, 64'ha74a7c1d046ab6e1, 64'hf1be3266e3a9d652, 64'h121f283e3d},{64'h1400000011900, 64'h170bc1100000000, 64'h7bcd9a61512cac00, 64'h34620ca8e2e8dd, 64'h5553f5d6e1d74418, 64'h15780042e8},{64'h8000040000c0, 64'h138206000004014, 64'hdccbba812c348f00, 64'hb86f96d8cdb7355d, 64'h20cc8b836d664de4, 64'h1aed994ddb},{64'h404000000000, 64'h116ac7400003008, 64'h9b4c4bc53c549700, 64'h26337be98926d3ce, 64'ha89e864bbe9b9f, 64'h16466a3770},{64'h20000, 64'h8737800000000000, 64'h29554de34081986d, 64'h6f0000007ff0f0de, 64'hcc46073202230ae4, 64'h7b8a60e01},{64'h6100000000040004, 64'h309bb56f62000014, 64'h9c61ae1c5c449651, 64'h592404376c51ed, 64'h8394e556b83d9648, 64'h1e9d},{64'h200000000000000, 64'h1734600000000c, 64'h9c537e2159000000, 64'hb44e464cdc658278, 64'h34bbdb92c66ed5aa, 64'h68004ab0},{64'h8000000, 64'h80b4000000001000, 64'hd6508e1b37deb275, 64'h837fc8dbe0006f4, 64'h448d51aa19190b, 64'hddf990c80},{64'h405008000100, 64'hf0f539b10800000c, 64'h98d3802d7a30984d, 64'hef13bb01b12c010f, 64'h9d322c06113bdae4, 64'h13d3},{64'h2000000100, 64'h117d00b18003000, 64'h70536d5970800000, 64'ha66c53b4e0800313, 64'he7b0c34c73dbd5, 64'h73d016180},{64'h400000000000, 64'h1ed5000000000010, 64'h3849989c48d09761, 64'h84a41cc708732bc, 64'h4d675bc5a5530fc9, 64'h84a5334d9},{64'h803010000000, 64'h3159829010000000, 64'h144992e37459e169, 64'h49331145152083fc, 64'h25048003f352435d, 64'h1c1a004308},{64'h3000000000, 64'h4579c5e000000010, 64'h4f8bab104c2ac1a2, 64'h6d3304fdb602727e, 64'he0dbb782090008bf, 64'hdc8286c9d},{64'h1000000000000, 64'h29a800000000000, 64'hda0ba3677b32488d, 64'haa6f46a8dc1b7348, 64'hb9381aa3e9abfbc9, 64'h4e09},{64'h2000000000, 64'ha800000000003004, 64'ha9d16ce179296cad, 64'h646c8581661603ef, 64'h912e947712001397, 64'haef8a1cbd},{64'hc050800, 64'h52c1000000004008, 64'h136d697c457271, 64'hcc37bb39b75bbd4c, 64'hed2277b160001ada, 64'hf8d004bbd},{64'h19406080040000, 64'h3000000000002000, 64'h42d1b4d706853871, 64'h4a143b457ca1426, 64'h20aee1ea61289035, 64'h10be141448},{64'h100c000000, 64'h3000000000004100, 64'h23129decb4d48a79, 64'h8c739dbd3808c4e4, 64'h2c0000059d6d90a5, 64'h50ea0b189},{64'h1800010000140, 64'h17acc0000000004, 64'h145d9e5c454200, 64'h735b840508a2369, 64'hb8ae8006bd289b7f, 64'h18e15d4efc},{64'h6000002000040182, 64'hc4cc4808000014, 64'hc6eb88285c3cb500, 64'h142b43786f709557, 64'haf85800428849086, 64'h81b0b1438},{64'h4000000004600000, 64'hc000000000000010, 64'ha289ab1cf8c89844, 64'ha54898b6000004e0, 64'hbf450006bc295bd0, 64'h1bd3792b38},{64'h201400000040000, 64'h2f17800000000080, 64'h6fc974105c589861, 64'h5d33000125eab5a4, 64'h1be6156ebb48f83, 64'h1946ccb7e0},{64'h440000000000, 64'h111000000004000, 64'h98ca95df5b360000, 64'hca01c9bc0726f556, 64'h856636137bd76cca, 64'h100f74704d},{64'h408000000000080, 64'h30d5c00910000000, 64'hd053bd6366489451, 64'h3c12c145818516e7, 64'h14075bbb33258f43, 64'h6f0a},{64'h500c00008010180, 64'hb159c9f018004000, 64'h9b6a262e5c469859, 64'h2b9b2993f5b499, 64'hed8255c3d1ad8a70, 64'h1b6ecc2b8d},{64'h61000000080, 64'h0, 64'hc08bae1506cde900, 64'h22ee5ac000000df, 64'hb094c6531c2817, 64'hbbb032c20},{64'h4004050000, 64'h3000000000000000, 64'h20ca6b2f14a09299, 64'h7a5936b526501b5a, 64'h503d00059c6e49c4, 64'hd70844dc6},{64'h8000100, 64'hc31626e00000000c, 64'hc8d69a04ac38987a, 64'h2b4e55295ad4a593, 64'h99bf0006fccadadb, 64'hb33122c95},{64'h301002000000800, 64'h1770000000000014, 64'hb00f4c59074c9541, 64'h6411022591f7ccda, 64'h69ce48929515844e, 64'h2d0004a11},{64'h601c20000040000, 64'h30b4443700005000, 64'h163e245c34b379, 64'h534c4142aec0eda, 64'h7c7f4ee4d9993b69, 64'h4476d2023},{64'hc01000000080, 64'h120800000000000, 64'h3b915ce09b29a000, 64'h122246b400000383, 64'ha6a5339f6e0d35, 64'haf8ef0000},{64'h100000c0, 64'h24d0000000001000, 64'ha98f9e10c15c8989, 64'hb01dd5700000037b, 64'h48a9000412ac16d2, 64'h84ee64a75},{64'h11406000030100, 64'hf117b80000000004, 64'h210b23264c24b885, 64'haf15ecfd1653f2a3, 64'hb904e19d4f4fd53c, 64'h9731f7074},{64'h10600000, 64'hb44a2000005100, 64'h10134e2af0dc9800, 64'h107db6d50ff318, 64'h5bc4fe3ee7d8c58, 64'h157db9bee1},{64'h200004000261800, 64'hbbd00000000014, 64'h7fd68614f755b800, 64'haf355deacddb8a8e, 64'h75386fb55e0005c6, 64'h157a1d5918},{64'h10400040, 64'h3000000000003000, 64'hc49badc8882d869, 64'h5f5d92b0501599, 64'h7b8741ee298530, 64'h1c54740640},{64'h509800000430000, 64'h5aab800000004380, 64'h7bcc3baa7c3c9049, 64'h5f59d4125860844c, 64'h39f7b9199d13a2, 64'h534f7c460},{64'h500000010600000, 64'h1008, 64'he04abd9f1806b800, 64'h6b928ac6214217, 64'ha92af106527d0db0, 64'h10a613145c},{64'h8000000, 64'h18504000000010, 64'h35497d5cd5dc9800, 64'h31935c6a0d74e5, 64'h748309d20c3c46a8, 64'h3289d01b2},{64'h1010a6000020000, 64'h6ad4ad2000000000, 64'h100c7ba14ba09899, 64'hf065db245155a206, 64'h205150b0c9357844, 64'h1b3041216b},{64'h4080050000, 64'h709b8aa000000018, 64'h6dd35e2d11a88d41, 64'h14e200f1b1710498, 64'hc585daa5140f077e, 64'hdc0001cf9},{64'h400000000000000, 64'h2b37800000000004, 64'h20d76a17613ac391, 64'h6a0ecc983b32746e, 64'h118671342a1a9bd4, 64'hf8a386f52},{64'h6000040002, 64'h12bbc5e000005000, 64'hb4b36d5c814894b1, 64'h6d3706d839db837f, 64'h814690a2da428fcd, 64'h7140f01e3},{64'h118005000001100, 64'h3091284000000000, 64'hd5be53ab8b161, 64'h3e05040137c0e8a3, 64'hf966782a04d68a4f, 64'h7137f62cd},{64'hc00000000000, 64'h8400000000004080, 64'h1b8b7a668748988a, 64'h6f6b8d91b23626f1, 64'h91bd9c1513705bd0, 64'h14742ef26},{64'h100000000000000, 64'h8149800000002000, 64'h1a91be1ab7aab064, 64'h59cb31ba86a6ea, 64'h34ae7036eaa9c000, 64'h16654d6065},{64'h400000008000000, 64'hf17aa82d0800100c, 64'h9c137ca8eb013802, 64'h282ef92cca3034e4, 64'hb92ed61e543e4dcb, 64'h181d1a2e16},{64'h2000010000, 64'h6b0000000000000, 64'h97e23575e7685, 64'h70624e293966e294, 64'h9cae327636e29676, 64'hd754f4a0c},{64'h400000020000, 64'hb137d8400000000c, 64'he8b73589c555104, 64'h196320e8a57793c2, 64'h70ee3196fde6d95f, 64'h1371e22cd7},{64'h14400106, 64'h1979a6c040000004, 64'h15b16caa5c3cb859, 64'h536df22729800119, 64'h49290510a2000afa, 64'h811001138},{64'h400000014000040, 64'h30e6800000006000, 64'hd6916510912cb881, 64'h78421417be2616db, 64'h38aee4e4de9e137a, 64'h18e77b2be5},{64'hc000000, 64'hc200000000002000, 64'h788f6c5d5826f452, 64'ha8225b70cd9e214c, 64'h70ce0002a4aecdc6, 64'h77c005cc6},{64'h4000010000, 64'hc6d4deae00000000, 64'hba3151158989b, 64'h1c614c24ae483108, 64'he0a9438638c2852f, 64'ha031c10a0},{64'h4000000040, 64'hd5a02000002000, 64'h3fcf9c9c98daaa00, 64'h616d6d859ff7827f, 64'h84a9f210a7daef, 64'h42f781c20},{64'h400405000000000, 64'hf68ae000006000, 64'h414e53132ac49300, 64'h55e0018c105652, 64'h49b0c523ef3b0cce, 64'h1ba72a31b1},{64'h6094441800, 64'h1b20800000000000, 64'h25957ded44823859, 64'haf92d58628efbbec, 64'h94fb9653ee000f46, 64'h9d89743b5},{64'h300002000000040, 64'h9b800000000000, 64'haf4b435967000000, 64'hbd000001652bd203, 64'h3a6601ef980536, 64'h1662b70000},{64'h1000000000, 64'hf000000000000008, 64'h75558de89405b80b, 64'h1464a778ea9de44d, 64'hbc3e12b2560013a6, 64'h778004293},{64'h4000000000, 64'h30e6ad0088005104, 64'h196285bccb561, 64'h436da90c6ab6d6da, 64'hc87900064a3543d6, 64'h42782e553},{64'h40000030100, 64'h3138da5590000000, 64'h168e2600bc51e103, 64'h5b0000006bec9647, 64'h6d6088620d196788, 64'h820865821},{64'h200005180000180, 64'h30d482a000000010, 64'h70488054665c8b89, 64'h66ebed78de9bc581, 64'h1c85ca039ed7d327, 64'hc38a00b56},{64'h100000010030080, 64'h30d4ad0000000000, 64'hc4cf9caa4a5c9871, 64'hcb34dafd88726515, 64'h139ed21eeb2c7ba, 64'hdc6ab5a60},{64'h400000000020000, 64'h107000000003004, 64'h150d4a9f38d6e000, 64'hfa4121503b6091c0, 64'h5129c0041cbe9072, 64'h11c5b942f8},{64'h1404100010000, 64'h6179c5e908003000, 64'h29922d565c02d871, 64'h6db16294dc75b318, 64'h1bf18d41342b585, 64'h1474b114e0},{64'h6000400014000000, 64'h7000000000002010, 64'h179aad26b2a049, 64'h9415f108d226f000, 64'h24a000205109320, 64'h14db825dd},{64'h4020000500c0, 64'h2716000000000010, 64'hb31586125c069879, 64'ha8000000d57096f9, 64'h41682bb383c29bd6, 64'h38776083b},{64'h803000000040, 64'h90800000000000, 64'h2d4b6b1f5c5e2000, 64'h3720cc190b56eb, 64'hcaa4c2c30ccb0c, 64'h138b1562a0},{64'h400000000000, 64'h277aa92000000010, 64'h991260d0d1509879, 64'h5d1c4975818e2654, 64'h6b38000655389322, 64'h18e2650654},{64'h460000000000, 64'h3138898000000000, 64'h1b127d6f048118b5, 64'h9d3706758ca04378, 64'hb593d9d2bbcb30b1, 64'hde9a842e1},{64'h300400000042800, 64'h30bbd00000002000, 64'h164a22d9c2aa91, 64'hc4633710db58c93a, 64'h6cee6126f54084e9, 64'h1ce57a2f46},{64'h2400000000001800, 64'h3026bc2000000014, 64'h2a915cd255409649, 64'h550aa00129d5fab8, 64'ha4ee620842584b0, 64'h1278ab13b4},{64'h8c020000, 64'h309bca3078004280, 64'hdc162e02dc011871, 64'h6fabf8b9be77007a, 64'hc41e83e338dc13c6, 64'h20d5bc5e7},{64'h8c00010000000, 64'h1ae0000000002000, 64'h135aaafbb098b1, 64'h79c70359d5134, 64'hacce6e6dbd1ad850, 64'h53c9b6141},{64'h4000005080000000, 64'h309b4c2000000010, 64'hc50501657d0b8a9, 64'h1cf3cca1b0b9d136, 64'h17c1304654000357, 64'h4e0321092},{64'h8010000, 64'h649ba2d410004014, 64'hdf936b985c5498a9, 64'h5c6c357dbc541282, 64'h6484d5f6fc000a0b, 64'h7ced01f5},{64'h300000000000000, 64'h7000000000001008, 64'he8deb0b357302, 64'h654a65949da5320b, 64'h9429653290000fb9, 64'h19576543dd},{64'h400000040000, 64'h3100800000000000, 64'h4b9174e4daa48b05, 64'h31462001b252e594, 64'hb2e613efca15ba, 64'h15f01f03e0},{64'h600000008000100, 64'h257aa92800000014, 64'haf76805e6c09a389, 64'h84e9d6cd537c0d5, 64'hed81d09000000e29, 64'he28e2607d},{64'h20040, 64'h3010, 64'h9408a42296ae7500, 64'h50000000ef6503ab, 64'hcd956b957200192a, 64'h3ecd635d3},{64'h1010000144, 64'h127b9a082440000, 64'h35758dc2b1800000, 64'hf371586d0d0b5295, 64'h101d8001e4b04835, 64'h1d8b64e04},{64'h60800000c000100, 64'h189abc2000005008, 64'h9cd48cd46c2dc041, 64'h5a0b7149af000075, 64'h7d376c1ebe001afa, 64'hf16740b7d},{64'h301000000011000, 64'h3000000000000000, 64'hcacea62f14c16099, 64'h64ec94dedc2d56, 64'he8ec00a3b48000, 64'h1963170000},{64'h1000000000, 64'h8000000000000000, 64'h34174a253105b87d, 64'h2a000000b4800412, 64'h84b49e32144a965d, 64'ha78d13c63},{64'h409802180000140, 64'h309bc5f600000000, 64'he0c451456b978a9, 64'heeb841504d8c3c5, 64'he400614aa5df8856, 64'h7100031a0},{64'h6400000000000000, 64'h1600000000005000, 64'h6fd3461550be42b9, 64'h9954a07d4f2a553e, 64'hc61c5bf03e0014f9, 64'ha050214f2},{64'h200104000c000000, 64'h2b37000000000014, 64'habcd8dd25c429691, 64'h98085ad15a0004df, 64'he6de00053f70ade9, 64'h1582bc2016},{64'h10410000, 64'h2800000000000000, 64'hc8c2e44013899, 64'hf155fb3b855ba42e, 64'h11685d712ec104b9, 64'hd4a183aec},{64'hc000040, 64'h1af5800000004008, 64'h38968a6a80389051, 64'hc2067b39668004e5, 64'h94e09a4280ae8a01, 64'h4bd400679},{64'h80000c000000, 64'hb0dc0000001000, 64'hc6c68f9b93000, 64'h659448715b8350, 64'h50c331464f5c4b88, 64'h132e1730cc},{64'h4001000004060000, 64'h20d5b143a8000014, 64'h418936016c4cb879, 64'h533bb510a59b492, 64'h5e6f800257add6a1, 64'hdee4a1df8},{64'h10061944, 64'h1200000000000004, 64'h277165e0f982b8b1, 64'h60487713b6d7aedb, 64'h12787d2c01f53c1, 64'hae93a2f50},{64'h400003004400000, 64'hf6810000005000, 64'h608e4c60cc000000, 64'h874e19e2be1d2306, 64'hd84349d30e2d8215, 64'h1657713282},{64'h418000000020040, 64'h30f5a42000000014, 64'hb2d5561c58ddb6a1, 64'hb82ba2e81ef0a6e1, 64'hbe5043ed702e89c2, 64'h16516030f8},{64'h404180000080, 64'h137c5d500000000, 64'hbed2826e8c000000, 64'hd6e15bec640000d7, 64'he8ddafb0d7ca07bd, 64'h5d0c96062},{64'h5004600100, 64'h709a2d0000006008, 64'h9c8c361ea034b3b9, 64'h8a709e7b260ba0a9, 64'hc45d0002bea297d6, 64'hdcd5b73d9},{64'h30002, 64'h4400000000000000, 64'h5075661f48ae9772, 64'h12a2848355c6fd, 64'h1b29652ba548508, 64'ha493c0000},{64'hc04000010000, 64'h3138304000000008, 64'hdb557b808c353891, 64'h2cb84d29e136f0, 64'he1bb3782cbdd84a4, 64'h165a066cba},{64'hc011000, 64'h1e00000000004000, 64'h504dbda69aa16061, 64'h1546300195674a10, 64'hddbd86f62a1bdae3, 64'h1bb5421ce2},{64'h100, 64'h30f6a6e000000014, 64'h974c80aca0b8b159, 64'h8842c8153900016b, 64'h5d3c8004f2220e2c, 64'h128a5e62b8},{64'h5010200000, 64'h1d17a00000000000, 64'h86929ae85c5c8961, 64'h344bb41a979614a1, 64'he93800d3e8581387, 64'h19a00d2624},{64'h300000000051000, 64'h62d4858000000010, 64'hc98f5d554c5dc041, 64'h3c0a44118cd048a4, 64'h6c1df194280f0288, 64'h1938000db9},{64'h1404008030000, 64'hf117804000001000, 64'h25d76a1c4c4cb80a, 64'hd26bf000296ac580, 64'h558642052ad096, 64'h13a7280c80},{64'h6014410000, 64'h1ed5242000004000, 64'h2b62351dcd861, 64'hb80abb2f93d04000, 64'hb8820f32d25484b5, 64'h55f2cb726},{64'h111000000000000, 64'hc, 64'h94d15a98dab9e000, 64'h5d64200190a53638, 64'hc0f1d0cb39c9dbf3, 64'h18e8b00032},{64'h8000014000000, 64'h68b4dea00000400c, 64'h9d62a1e5c422291, 64'hf76396fd4f827202, 64'h883d8dd3e0cc810, 64'h4ddb90734},{64'h61800, 64'h317a856000004280, 64'h168c269051c279, 64'he5618795b0ea5800, 64'h8d8618d378635861, 64'h1949cd606},{64'h800000030000, 64'h138bdaa08001000, 64'h6a50649cb0000000, 64'h630000015a53d374, 64'hec4b8005a17d04b1, 64'h1586fb2c8b},{64'h300004000000000, 64'hf0b4800000000000, 64'h6911aaad70b20203, 64'h2806740f99d59a, 64'hebecb576704fbc, 64'h10c4200000},{64'h2000000100, 64'h5359c84000006014, 64'h7dd6705a6c3ee0a1, 64'hf7338000ce1fe25d, 64'h610c241338904a05, 64'h15f5f803f8},{64'h8003008000000, 64'hf6800000000000, 64'h61cbab24ea5e2900, 64'had229c9c689871a2, 64'h10bdbdb382b4b8c, 64'h15c2d55aa0},{64'h1400010261000, 64'h557ac5f6a0007180, 64'h4f133604ec051849, 64'h8c001b5392dc4a0d, 64'h34000005732dc5b0, 64'h6b64a96e2},{64'h1420000000000, 64'h1e00000000004000, 64'hdb0b8e204c02f851, 64'hbe30e60dbc0be3a4, 64'he8ca8a05839eab04, 64'h5b7766f0d},{64'h1000000000, 64'h4558c82000003000, 64'hb4e157a59809b, 64'hed2149d885196380, 64'h4d980004eecc0c3c, 64'hbedc14a0c},{64'h0, 64'h6800000000000004, 64'hbecc5be6a75aa994, 64'h93652be895007254, 64'h5d0a2fc19c24c670, 64'hb0408599c},{64'h5008000180, 64'hda9ac5f07000400c, 64'h1f5258586c50b6bc, 64'hbbdf7979b207d413, 64'hcb314b2cc000955, 64'h68e725f9e},{64'h100c000000, 64'h17a800000000000, 64'h7cc6b974c266200, 64'h382bfd39a2038278, 64'hbc100cd2ca335454, 64'hae800177e},{64'h10200000, 64'h3158bda040003000, 64'hb24eb0ae462c93a1, 64'hdd03f59baf244596, 64'hdb0000238911bb0, 64'h4b7602389},{64'hc00000010000, 64'hc501800000000000, 64'h804f5d5517268cb5, 64'h62a69509ce46f1, 64'h8d2a026eddecd28, 64'h728e46ce8},{64'h119002000000000, 64'h8121000000000000, 64'h9e0bbb60c9d5287a, 64'h6542096d0b2784de, 64'hb084cb7e099958ae, 64'h960004bc4},{64'hc00000000140, 64'h30b4284000001110, 64'h2ad59de9203c91b1, 64'h8637e6189e0ab1c5, 64'h40df0d04f36f8b01, 64'h139e5eccb3},{64'h428403008000180, 64'h5f7ab56000000000, 64'h529236214044b361, 64'h144378b98ca2e371, 64'h998a586a630019a6, 64'hf884b0965},{64'h86, 64'ha4862000000000, 64'h9d2bbe268a829800, 64'hae436b3c3f2cf209, 64'hfaab60fc6b8559, 64'h193e1b0fc0},{64'h2001060000000000, 64'h3117c06000002014, 64'h136d52c9288ea1, 64'h16c42165db81c4, 64'h4fbe1090fb2ae8b8, 64'h4c4b72bbb},{64'h1000000011000, 64'h120a800000005000, 64'h9950b62766b0b891, 64'hac2442b082569974, 64'h885d8c116db716e0, 64'h1b8e6663a4},{64'h5090061800, 64'h309bce2a00000100, 64'h1a8f2c2c462c9269, 64'h2797532585721bec, 64'h11006b4401ad5c7, 64'h18ef7fa040},{64'h3000000044, 64'h5000000004014, 64'ha7edbbd9674c9800, 64'hbc1602bd861a337f, 64'h516a0cf16033c19d, 64'h64eaa175b},{64'h0, 64'hf6d00000000000, 64'ha7ce9c969646a100, 64'hba6198710e0002c6, 64'h10ae8a8174000f90, 64'hc22a01506},{64'h500402010600000, 64'h171726e000000000, 64'h4c13852cc0288d41, 64'h301438676592f2c6, 64'hd1b2ebc377b044bd, 64'h1670b42ba2},{64'h2000000000, 64'hc2b4800000003000, 64'h1d51adecac21a0a3, 64'h3b47654882152338, 64'h587f0563fe410e16, 64'h104763f01},{64'h1000000010000, 64'h24d5d66a15825100, 64'h384f6500ec5c8989, 64'h172be414ce72720c, 64'hc50c4000df854afa, 64'ha15f8aba7},{64'h4008000040, 64'ha80000000500c, 64'h8cf5c677b415200, 64'hd5abe4406b84389, 64'hdc1180072408c444, 64'h128c245ab9},{64'h401460000000040, 64'h309bbd8000000008, 64'hf4b2e224a4c8ea9, 64'h5a2d0169b693d16d, 64'hd406f784e12de46c, 64'h5a8002c52},{64'h40000500c0, 64'hb44e2000002000, 64'h3192ae1b40dc9800, 64'h970ca319afe76307, 64'h21bd4941280201e5, 64'he9e511dc0},{64'h400000000030000, 64'h3179bd6e68005100, 64'h154846ac0a3891, 64'h9d13a800856136b4, 64'h743261e661e15030, 64'h1945c193a8},{64'h300000000000080, 64'h200000000000000, 64'h960fb61736c552ac, 64'h7b47a2491e892255, 64'h17e6726555ed301, 64'ha72590000},{64'h100000000000140, 64'h5359d24000000010, 64'ha0d80808c3c91b9, 64'h21050629948214a7, 64'h1c1c292cdca8c50, 64'h84b181610},{64'h508003008000100, 64'h3158ce0000000000, 64'h79544bd05c489769, 64'h7169d634c6ab404f, 64'h3081420ee2001a2f, 64'hf33712cfb},{64'h201420010000000, 64'hb0b1800000003018, 64'h94ce4c665a5c88a9, 64'h7b3cb155227671c8, 64'h51b065431b472723, 64'h1664575619},{64'h4000000, 64'h4600000000000010, 64'h50099e1776da028d, 64'h4134b994d080042c, 64'h750165c082001090, 64'ha0a9d5f7a},{64'h2014040000, 64'h30b4c5d310003000, 64'he056806e5401b8a1, 64'h7a281b48ced604f1, 64'hc1bcb6570803532f, 64'h1385485a6a},{64'h1060008000000, 64'h4200000000000000, 64'h4a977ba6b531b1aa, 64'h30d5c0dfcad15a, 64'h20691884836fab80, 64'h958001a46},{64'h500001010c, 64'h668b800000000008, 64'h34752d94662c8d81, 64'hf934a001175a530f, 64'h350dacc11a23056d, 64'hb3ecc6512},{64'h8000000000c0, 64'h159352000000000, 64'h6fcb7b9910800000, 64'h8410600167d9d0fd, 64'h600840fd408df8, 64'h848c00000},{64'h800014040000, 64'h1800000000003000, 64'h218d94615ba1e149, 64'ha030f8f85f51ad3c, 64'h1d952026f98091f2, 64'h5bf285402},{64'h1000000080000c0, 64'hbbce0f68000000, 64'h338ab4589c000000, 64'hf724561867186183, 64'h405dde60127996e5, 64'h880000124},{64'h25300000000, 64'h9759bda000004100, 64'ha0018e286ba88e41, 64'hced0497d5530a270, 64'h81859600d788249c, 64'h44cae165},{64'h100002000000100, 64'h3000000000000000, 64'h58d79c9766aaac0d, 64'h5f161190b18640fb, 64'h416a5f3020000ded, 64'ha103d07a0},{64'h2014c0000040000, 64'h70e5d66a4800000c, 64'h1440626c5cd803, 64'hb01602581c61cbd0, 64'hc05449719b576f40, 64'h1661e93092},{64'h4008000000, 64'h34000000001000, 64'h6d0d9e22b95a0900, 64'h459d0559632b261, 64'h1c1b65376055bb5, 64'hb25bb2000},{64'h10600000, 64'h2937800000002004, 64'hac0c6e13774540a9, 64'hb062b8eeafab020a, 64'hb4000002589e4962, 64'h3b5604333},{64'ha000000008000000, 64'h7141244000000010, 64'h5e158decb0b89079, 64'hd02bf340bc1a820e, 64'h7a3d29a0f4a690bc, 64'h841bd2599},{64'h500800000010100, 64'h2ef6b9800000000c, 64'h12c9ae2259d8a8a1, 64'hc232e1e006c78157, 64'h3068677f2586c261, 64'he080070b1},{64'h4000000014010000, 64'h3159800000000010, 64'h8945e5c5c8b81, 64'h4295a7bc5ae35c, 64'hfb2a8ae2163c0858, 64'h13b8af0970},{64'h4280011800, 64'h5200000000000008, 64'h42ce7c10c0549669, 64'habb7e00085c6593a, 64'hdd9c4388428d74, 64'hcc8e13830},{64'h1000000080000c0, 64'h3161000000000010, 64'h2b0f4dda87309891, 64'h213b2b990802429, 64'hed0f47b4e4984570, 64'h1c3cad3731},{64'h1114000000, 64'hb158b56000004198, 64'hc60e782e54c0b3a1, 64'h7b959411afa1c652, 64'h81b021e3e6000b35, 64'h133659e3bd},{64'hc04000000080, 64'h3000000000000004, 64'h63557357465ae099, 64'h396e233c67b10051, 64'h9888038053440814, 64'h2137},{64'h10000000508c0, 64'h71205c2b10002000, 64'h85116e264a308fa9, 64'h146f60018658dd6b, 64'h89b412219f951b8e, 64'hf34001ca4},{64'h8004000000000, 64'h178a84f08005100, 64'h25d260d646800000, 64'hb46de259a9b786a6, 64'h602be54968de05d4, 64'h1504e5a822},{64'hc000080, 64'h2ca0800000001010, 64'h71179adf2ab891a1, 64'h6b345de9978004f3, 64'h5fc13033f01acfc0, 64'ha0c0f1698},{64'h24000020000519c0, 64'h4117cc4000000018, 64'h9cd46e1c685cf862, 64'hd265c968a9561b39, 64'h4e2b601402001bd4, 64'h100a753f1b},{64'h11000000c000100, 64'h110800000000000, 64'h2b779a5a87489800, 64'h2a2e10a90a02464f, 64'h869588c36000120, 64'h1210000489},{64'h1400000000000, 64'h26b4000000004000, 64'hea0545854b889, 64'hef0baa4d498ef1de, 64'hd85b0000472362e8, 64'h127546a82},{64'h218000014000040, 64'h68c5800000000010, 64'h2b558d924540b299, 64'h20b52504a39f37f, 64'hb884cc0800000425, 64'h6410916b2},{64'h14c0080000100, 64'h70bb800000000000, 64'hd7498e266a2098a9, 64'h2ac28e09c13ae18d, 64'h5dce368011253507, 64'h67a173f08},{64'h800000000040, 64'hb08080000000000c, 64'h9d556b277a264b02, 64'hd43a82753a89d19d, 64'hf96a000013c2d105, 64'h11f2ab2218},{64'h110c00000042800, 64'h7159bc4000000000, 64'h63c82ae85bc49262, 64'h9950557c4963db14, 64'h74b070bda9a6593a, 64'hc5990650c},{64'h2000000140400c0, 64'h117866000000000, 64'hb4905aac545ca900, 64'h763156f410cb0439, 64'ha4b277a6f40004bb, 64'hde9a92c97},{64'h4000000, 64'hb1542080002010, 64'h67084cdb175c9800, 64'h88161410db00037e, 64'hec8118837eb3d679, 64'hf4ea95996},{64'h30000, 64'h516800000000000, 64'hf4c1d7b2e819b, 64'ha559c1d19652c000, 64'hf43980053aa954ea, 64'h1c26b159ca},{64'h300005118000002, 64'h2290544000000010, 64'h41b36614b9389079, 64'h2cccb9cc68273561, 64'h93d64d00000020d, 64'he11a753b7},{64'h40000c0, 64'h140800000002000, 64'h4c084ae6da800000, 64'h4c1a1000261302f1, 64'h425905260414cc0, 64'h844de37b7},{64'h100c000000, 64'h2800000000004008, 64'h620d4beaebae008b, 64'hce099621561682d0, 64'hcc000005c24fd0de, 64'h95daf0993},{64'h500400000040080, 64'h3179a44000003000, 64'h38557da25c017875, 64'ha4e0994d2d6635d, 64'hed6663f4ef8fc85d, 64'h57e702ca4},{64'h400008000000, 64'hf6800000003000, 64'h244a5d533946e000, 64'h873771a04886847c, 64'h568873899b1390, 64'he063f4560},{64'h18000144000c0, 64'h2359de8c08001010, 64'hc8d0782c54a8d869, 64'ha547d2ba39800645, 64'hd053074405d80530, 64'h56f2a10f1},{64'h9400000040000, 64'hf0800000003000, 64'h434ba3591826e200, 64'he42ee4e4c343919e, 64'h10f760bcd0e01c8, 64'h82d0e2ee0},{64'h800000610000, 64'h160800000000000, 64'h40a9caf14c1f500, 64'h1f073c4667f7b6d0, 64'h3286422107c080, 64'h32af35e60},{64'h101000000050000, 64'h9517800000000018, 64'h3215b010d6409749, 64'hce16800c324c85a4, 64'h4c916cc02100dbc2, 64'h1ba00007bb},{64'h10020000000c0, 64'h3137deb210000000, 64'h5966ae080c498b1, 64'h993f0001bf3616a7, 64'h5c0b0625997105a5, 64'h1bf8621310},{64'hc01010000000, 64'h16d4c82000000000, 64'had94aa1f113098b9, 64'h102b000832cf20c, 64'h19957770927cfc6, 64'hb210013e0},{64'h400000041000, 64'h70f5442000005000, 64'h15be289b349841, 64'h385f60e0aff2eb12, 64'h283e18a4031f17d8, 64'hb0675df66},{64'h10a1000600000, 64'h138800000002000, 64'h870bb360a930af00, 64'h494370aaa4a9e292, 64'h10f1f45351ea125, 64'h12cf05400},{64'h8041800, 64'h90000000000004, 64'haae2ed6523600, 64'hbd0bb6d83c6939df, 64'hdd0c9f44ee6f5381, 64'h4aa186a99},{64'h300040000010000, 64'h80800000000000, 64'hbdc96b1f38ae0e00, 64'h9e110bdc4a55f10e, 64'h91d06172133230b8, 64'hb208913c5},{64'hc010100, 64'h179b45010000008, 64'haad2b25155a89100, 64'h844411edc140013b, 64'ha1ce63e5a82103d8, 64'h11408442f8},{64'h500000008040040, 64'h56d0000000000000, 64'h8acf4c6059bae341, 64'h603a92f8017274eb, 64'h3dd8b0c081c5f0, 64'h1c036747de},{64'h0, 64'h1174e00ab421100, 64'h34d77e1095800000, 64'he33c6b0469ac1352, 64'hb0c80006f8640f59, 64'hc5d90b7a7},{64'h400010000140, 64'h9759de9288002018, 64'h6e0e26156030af81, 64'h3b6e3b5c1d80031b, 64'hddaac6f586d6b8, 64'h169e173cd0},{64'h1800000030102, 64'h3148800000000014, 64'h6ff06cd971249879, 64'hb53a28482782429, 64'h88058004a9d7967c, 64'h1c20a21cb2},{64'h2184000000, 64'h116484000000010, 64'hdec99aeaf4000000, 64'ha5d9d1a83a46b118, 64'h4046b6e11a0014ee, 64'h3637c2839},{64'h4014010000, 64'hf000000000000000, 64'h58576a596756680a, 64'h396f56d939d04208, 64'h28b020a38400035d, 64'h989053858},{64'h4000030040, 64'hd5a6b6aa020000, 64'hcb8c8ddd31000000, 64'h4259c00026706261, 64'h856706120b908696, 64'ha032e5901},{64'h8610000, 64'h22d5800000000010, 64'h4b09add8a9011879, 64'h2e217b936750a2d1, 64'hb9380ee1ac4b86b1, 64'h6b12d4854},{64'h400000000000000, 64'h9b858000000000, 64'hb8f5c5c8855a200, 64'h8a4e45c0b370565e, 64'hbc5b66e2c2228b08, 64'h19814e47e0},{64'h3000000000, 64'h30bbc5ea08001110, 64'h568e4c2d5449a099, 64'h3f14c58592961212, 64'ha91f8000e843043e, 64'h11fe2d95dc},{64'h1000000000, 64'h116482e00004000, 64'h1213bd5741588f00, 64'h106165d9858f71ee, 64'hb83a5e362078c537, 64'h67c491ca2},{64'h1400000041000, 64'h629bdaaf68001000, 64'h122d02ac4d6071, 64'h466f8de84ec39800, 64'h3cbbada6171193c0, 64'h8767a5b49},{64'h100004000000144, 64'h1b1780000000000c, 64'h4305a653030b851, 64'h766f008857a432bf, 64'h1032cb10440014cf, 64'h58a435e79},{64'h300000018050080, 64'h137000000000010, 64'h57c8a36a95ca2100, 64'h3212f4345850d59d, 64'h4f69d641c40c91a8, 64'h11b9643d3b},{64'h404008000000, 64'h11780000000000c, 64'h1993755376c08800, 64'h202d198ec9f40fa, 64'h80ed87e38b1f8c45, 64'h1bfe2002f8},{64'h860000050040, 64'h5979800000004000, 64'h1b8db3d3558638a1, 64'h705a1394966fb20d, 64'hc0000002ef592728, 64'h158d081ca1},{64'h800004040000, 64'h150800000000000, 64'hdb4bbc60a9a49800, 64'h75f7e70686d2734, 64'h4cc572b0f9849963, 64'ha52b143cb},{64'h80, 64'hc281000000000000, 64'h9d96bcdb18552b53, 64'h790f21a43486a293, 64'h890c1da541950ff8, 64'h3106b3721},{64'h1000000100, 64'h309ad26b44a25000, 64'h2217789900055869, 64'h882c68fd1f853311, 64'h212418a314000dec, 64'hd7c542829},{64'h1002000000000, 64'h189ab9a000000000, 64'hbe12506f104c9459, 64'h1082b939af80f6, 64'h491d447f7504f4, 64'h13aa501240},{64'h6600000004040140, 64'h5f7ac81608000008, 64'h2c944a14564cd869, 64'h650f7d8034760123, 64'ha256c526ca144427, 64'h290b35ad8},{64'h1000000000000, 64'h9b800000000004, 64'hdc487b664ab89100, 64'hcb6e2948db166276, 64'hf0b28cb6c16f5164, 64'h1b927c7019},{64'h800000000100, 64'h31680000000000c, 64'h6ec99aef2432d57d, 64'hbb376650ddaac19f, 64'h5cf1000321789be5, 64'hde1e23d98},{64'h404000030000, 64'h110c8225d020000, 64'h120c4bef3402b800, 64'he45afde90dc036a6, 64'h24510ca3777900fd, 64'h20bf17e1},{64'h10c00140, 64'h10bbc5ea4b001000, 64'h1ac19e1a5c58d8a9, 64'h6b0072d3b7283191, 64'ha9420280c60a0468, 64'h1c276a145d},{64'h400460014000000, 64'h18b4bdb008000000, 64'ha62f113898a9, 64'ha73f1b30cb89f000, 64'ha43176911b9d64fa, 64'h1be5c1372d},{64'h1005080000000, 64'h2ad5800000000000, 64'h20538e134c055881, 64'hc2a80c1d210812c3, 64'ha40000013fb3900d, 64'h1652e965cb},{64'h3010000000, 64'h177ad06000002000, 64'hf40452c2a6049, 64'h5007135885a7b4f6, 64'h7c85af5040001216, 64'hb4d005ea0},{64'h80000000, 64'h30d54c2000004000, 64'he5e2b1b512261, 64'hd6c367e139306000, 64'h78828c94e0324974, 64'h785074363},{64'h0, 64'h70f680000000408c, 64'h208c5a553951c20d, 64'h1b15a0011708264e, 64'h7d9509f2ba2b4b0e, 64'h4af30aed2},{64'h500806000000100, 64'hb127b577a8000000, 64'hc2ccb0685c44d803, 64'h764407e0b0cde5ef, 64'hd90bcad2194150bd, 64'h81af620ab},{64'h400003000000000, 64'h44b4dc0000000004, 64'ha74fae11554a788b, 64'h1d65c2fd85e9d6f8, 64'h6d1f72a17ec75887, 64'hc829b21da},{64'h718004114010000, 64'hf117deab4d820018, 64'h60cd36246c38b341, 64'h7797d90dbe4b06f0, 64'hc4c5edab0627c305, 64'h13d6446512},{64'h18041140, 64'h161000000000000, 64'h388e7dd330aea000, 64'ha03c74b960f789a7, 64'hbd6aaba540b54972, 64'h15010620e3},{64'h100000000040000, 64'hf138000000002000, 64'he1cc6bd2b5391105, 64'h2354602c1dd0d816, 64'h38b244708e0383f0, 64'h11bea30480},{64'h300044014000000, 64'h30f5b9b000000004, 64'ha8e12594c96b9, 64'h1453bc5072b41130, 64'hcedf140fd41e05f, 64'h1a1099441c},{64'h4000000, 64'h9b502000000008, 64'h26516ceab4000000, 64'ha1cb8286289918a, 64'h4824000656470386, 64'h240c6211c},{64'h418000000000180, 64'h709a3117ada85388, 64'hae0e585e6c449379, 64'hb87391855c313209, 64'h650561ec24cc030a, 64'h82d31da78},{64'h400003000000000, 64'h2600000000002000, 64'h320fae291badc181, 64'h7e2fc32539000192, 64'h2430d644ef590ed5, 64'hdf6404ee2},{64'h300000014020000, 64'h24d02c2f02444080, 64'h9d53bda85c28b889, 64'hdb4e176d1fc8a114, 64'h12463e124925251, 64'h96c89ac90},{64'hc100865000000000, 64'h66e0800000000010, 64'h20152d9ed85db889, 64'h64f22003b2466c0, 64'hfe4966115f752457, 64'h13af3005f8},{64'h1804114010000, 64'h3179d82000000000, 64'h126e131c50d8a9, 64'h6594d169b053c05c, 64'h6c296530e95951ff, 64'h2d82f6e41},{64'h180000c000140, 64'h9b282000004080, 64'h41089adf5101b800, 64'he737bb9d7583b1ef, 64'h24848003c7654f12, 64'h24f72cf94},{64'h4008000000, 64'hf100000000001000, 64'h14ae177644930b, 64'hca5b10016809d000, 64'h786509e3c5b3c234, 64'hde4c95522},{64'h440010000000, 64'h3000, 64'hc5cc4c5756bd5400, 64'h510451498ba200a4, 64'hb110800195d57030, 64'h272c7091},{64'h300004000020000, 64'h30b0800000001000, 64'hb5c9be271b560c4d, 64'h3655066031ed7598, 64'h54246755c0d8194, 64'h364676fb7},{64'h30100, 64'h1b17800000000008, 64'h1d1575ed202e6149, 64'h80e80004fc380cd, 64'h31970520a41cd673, 64'h174800387b},{64'h6000000000040000, 64'h70e6800000000004, 64'h1b127de0b0322245, 64'h6d5720017deb92c0, 64'ha66580057232c811, 64'hb106d2d3b},{64'h44, 64'h30f626e00000400c, 64'h42f2756c440a1889, 64'h1b1bc8e11c08d4f7, 64'h10ba7320a230106, 64'ha56732190},{64'h1c050086, 64'he891344000004018, 64'hcc757e22c0ba4099, 64'h310f362034d884e5, 64'h50000000a84c5951, 64'h35d310c51},{64'h301400000000044, 64'h159c00000004000, 64'h86ef4c5647000000, 64'h5f09617c8215245d, 64'h4cb15f5315caa258, 64'h2a5534405},{64'h1460010c, 64'h138ca01a0000000, 64'h1ee9aad4d1000000, 64'h8c1095de469a95f1, 64'hf4599bd6542cc83c, 64'hb408e2d06},{64'h3008000000, 64'h1407000000004080, 64'h430bab6914b08f41, 64'he917f32c20800196, 64'h5220001627a4c85, 64'h59f2fbd21},{64'h200004000000000, 64'h30c0b84000000004, 64'hbd945e1ea8cc96b9, 64'ha354028d172f6307, 64'h1858c710e200065c, 64'he98f04894},{64'h1804114071800, 64'hb0e6deb38c840000, 64'h8261690a0b8a1, 64'ha0b77000ddd0e800, 64'hd85404a42fb56dde, 64'h612361848},{64'hc700005180200080, 64'h3000000000000010, 64'h9ecc3e106524ab69, 64'h88849a8f8a341017, 64'hfe51703684b54f27, 64'h128abd0932},{64'h1406000000000, 64'h140000000001010, 64'h75556b9e9c5d1800, 64'h2b6292118920a2cc, 64'h18b300005152c46f, 64'h1a17866d5e},{64'h400001008600000, 64'h1751000000000000, 64'h85179e18fb468049, 64'h1b4154730d8000c2, 64'h25b4c8242e4248e6, 64'h15c9051044},{64'h20000000c050102, 64'hf080d86000000000, 64'hae2b4be2ea288d15, 64'hc50c3bd521441103, 64'hb90cf2d663cb57a9, 64'h2104138a6},{64'h400002014600000, 64'h1e00000000000004, 64'h6fd54a14b8c09369, 64'hbb1ad5fadf9bb193, 64'h2d7ae5b0000013bd, 64'h13aa744e72},{64'h20100100c000000, 64'hb0000000000000, 64'h1d4ae12d4523700, 64'h9f3b727c56807115, 64'h4d3b483193001254, 64'h1a98ae106d},{64'h6500000010000184, 64'h137a800000000004, 64'h1daa336259a0cba1, 64'hf015b6ed3cdbf105, 64'h1e4fc5b5ec42d7b0, 64'he010c6619},{64'h200000000010140, 64'hd0000000000010, 64'hc74f8a6b34389000, 64'ha2544000b371d617, 64'h6f3e73f536cfd4da, 64'h5ed1},{64'h610000400800014e, 64'h1e00000000000018, 64'hdf3525dc6844d269, 64'hcf5cf6f55580053b, 64'hfa84d956f42798ee, 64'h1765bc5376},{64'h100000000000100, 64'hf0800000000000, 64'h9c896cdc4c468200, 64'h372ca9e18c1666f1, 64'h244f42d05a0dc654, 64'h13d2504e65},{64'h200000010000040, 64'h117b9aab800000c, 64'h134a24ba8e8000, 64'h25d11c3f0470a5, 64'hc110ef00000003e8, 64'h15787f659b},{64'h3010a6000000004, 64'h5b17000000001000, 64'h70a0462904ccb559, 64'hc3386289670a25af, 64'h3833ca201d11e3f5, 64'h167ce61cc4},{64'h4051804, 64'h2540800000004000, 64'hcbb36d52552cb889, 64'h59d12072ee98e9, 64'h686309a090318000, 64'h4cc0018c2},{64'h50000218000018e, 64'h1e00000000004080, 64'h316a3b1666b8b351, 64'h6fad23195ccc6133, 64'h42440020c3c8865, 64'h63562ad25},{64'h4030000, 64'h159800000000000, 64'h94ca5c9cf1000000, 64'h854374c51c75a11b, 64'hed2427c70a1ed773, 64'h1768480901},{64'h401820000000000, 64'hf0f5a93300007014, 64'hb38eac5b7c20f061, 64'h59ce0dc1b6c12a, 64'h54b25532c915298c, 64'h1206cf1132},{64'h2001000000000000, 64'h995e4d00000000, 64'hae53ad164b000000, 64'h281664ad5c92b11a, 64'h8640a281254ac46a, 64'h408002a78},{64'h80000000010a, 64'h237a48400000000c, 64'hd8337d6d00a08c69, 64'h3d26f0de9a5101, 64'hd4dec2f1670bc040, 64'h19a8082d1c},{64'h1180000080, 64'h1720800000004014, 64'hd8104e275a348f41, 64'hdbdadf8f70be197, 64'ha5c00017e2e0f4d, 64'h17f7f6e51},{64'h2200004000000000, 64'hf6000000003000, 64'hc2ceae2774c89400, 64'h3c0aa0f42b2a565c, 64'h1ee9c3d65c158f14, 64'h117ea03a74},{64'h400000000c000000, 64'hec00000000000004, 64'h86d54e1b19be5475, 64'hf309586d0e2d9294, 64'hdb6c8481511b0361, 64'hb11611858},{64'h1000000080, 64'h2179800000000010, 64'hd8c6d691c26c879, 64'h7c64a2981b0004f9, 64'h9d31000685cb16ae, 64'h53a7d0d92},{64'h4000000040, 64'h2e0000000000000c, 64'h1bd1625135be42a1, 64'h7b436210378b02cd, 64'h14000001041bc1b5, 64'heb48570d2},{64'h201000000030000, 64'h19384000000000, 64'h4311ae1335d1f700, 64'h7c0000010cef5082, 64'hc8415c50a542620b, 64'hd790d6fad},{64'h1060008000000, 64'h1351000000005000, 64'h37115a9a80da00b9, 64'hf95ebbe57c8004e8, 64'h293b800197cb7452, 64'h36d0a4dc4},{64'h500000000000080, 64'h7148ce2010004000, 64'h27c9baeca0c09861, 64'hac01ad9c4f8ac37f, 64'h139dda106768068, 64'h139f4201ae},{64'h5004040000, 64'h1f58b8170d023008, 64'ha2cb9e20a924b869, 64'hb13fbd8c468b37e, 64'h2441cf33a6749955, 64'h574956a74},{64'h2010a00000, 64'h2e1b4c4000000018, 64'haa8f4ba2d02cd8a9, 64'h770bf12f4dad52c2, 64'h84b22d42985dd7b5, 64'h18f34220b5},{64'hc01010400000, 64'h3080502000000000, 64'h6d0dbd5ec8add649, 64'h7a655a8b67afb63b, 64'h84deafc67f1854df, 64'h15ba4a5f81},{64'h401400000000000, 64'h30f5862000000000, 64'ha80aab688132e049, 64'h4e2cc13d3c25b2b4, 64'hc9226f7163138278, 64'h1508b25ee2},{64'h201000018e00140, 64'h5b17ce0b48000000, 64'h1f92b069505ce851, 64'h147a825d1a95ed, 64'h9966770e39dc3f0, 64'h1398bb1747},{64'h300000000020000, 64'h200000000000000, 64'h33cbae28a4b50fbc, 64'h7365422423f2e144, 64'h31784e64e644044a, 64'h16c72f1129},{64'h20000000c040000, 64'h92d0d80000000004, 64'h880fbe1cb8c153ac, 64'hc6387abd8a4a2c12, 64'h18876213a8249070, 64'h16c0861cd2},{64'h8000008040000, 64'hb0b4c40300000000, 64'hbce7e2f66a27885, 64'h340910e10542f59e, 64'h6349aac80d16e0, 64'h1688390720},{64'h140, 64'h3117dea000004080, 64'h99aac4401d881, 64'h332d3ccdada420c3, 64'h31768cc198001adb, 64'h15cd07e143},{64'h300400000000000, 64'h44e5b56000000000, 64'h19154c10c029865, 64'h8f3b685d0b9372c8, 64'h1d24c904f97c1c2c, 64'hb28000000},{64'h40, 64'h30bba92000000010, 64'h4ad6aa26fa448d91, 64'h500a0201c1c8012b, 64'h3879b33666000830, 64'h83b081172},{64'h200003000000100, 64'h159ca3702c21000, 64'ha4cd4ba0c4000000, 64'h3505e17495e9300f, 64'hf040ed0000001147, 64'h4773505ea},{64'h400800000010000, 64'ha32100000000000c, 64'h428d5e264c54974a, 64'h12e3b8deded011, 64'h602dc9a05f78c4d0, 64'h4c10b66b2},{64'h0, 64'h106800000001000, 64'h179a5125d5e200, 64'h3d0aca805ff0c536, 64'h2b240480001970, 64'h1bfe9c07a9},{64'h1000000000000, 64'hf0e5a6cd58000000, 64'h8710a8e4c1454104, 64'h6705a19c3602d54b, 64'hb81700013d7d1450, 64'h198b166620},{64'h1404180000000, 64'hc338b17418002018, 64'he8c84aa06c48b5bb, 64'h6ccf89956cfa3000, 64'h53ba905bea41bc, 64'hb14014e70},{64'h41000000c0, 64'h2ec0800000000004, 64'h1d12982c44b48fa9, 64'h2cb840003a1c006d, 64'h5042ae61621d0007, 64'h3800014f6},{64'h40080, 64'hb081302000000004, 64'h9f155ca8fbb49803, 64'h292f7e016777c0df, 64'h8148004f8951c00, 64'h1b602810b1},{64'h1000000000, 64'haac4000002180, 64'h3dcc4c6089b9f700, 64'h724e0375bfb596fe, 64'he47c0b90e42e4e2c, 64'h2150d9f02},{64'h8640000, 64'hf0f5c5cd58001000, 64'h34abb295b065804, 64'h7b5159de6347b262, 64'h116c8c4090b64240, 64'h13ad322153},{64'h4001060018200000, 64'h5ed5dc2000000014, 64'h5956325c58449561, 64'h492630365b16516a, 64'hb730000f776a5b1, 64'h1c0ed3091d},{64'h600002000000146, 64'h7000000000004080, 64'ha2f58de16a249861, 64'hc13821995586659d, 64'ha0a9da53a7b5084d, 64'h167d0cdaa5},{64'h300001014000104, 64'h7159800000000000, 64'h58716c9f40289859, 64'h77167ca16732a573, 64'hcda16775f8c10bbe, 64'h1698005a69},{64'h10410000, 64'he000000000000c, 64'hb3937d5ab8a28a00, 64'h3d36f76875f4f0, 64'h857e6d34b85757b8, 64'h169b89495a},{64'h301000000000000, 64'hf0b1406000002000, 64'hdf09ae1176d9c103, 64'h244ee910b3644174, 64'h117be441710905d0, 64'h150c240fee},{64'h800000000000, 64'h321286000003000, 64'hb24f4c577c4db5b4, 64'h4d5a013444ad0498, 64'h28e14354ef0d46e8, 64'h3fd0c4424},{64'h88000100, 64'hb0f6ce3410003000, 64'hebeb82657aa8980d, 64'h7391390505241437, 64'h602c0004822ec886, 64'h197e211741},{64'hc000000, 64'hc5800000000008, 64'h850f5626eaa68100, 64'h2241f85cea61e572, 64'h701ca1e432088f80, 64'h1680005b18},{64'h1403000040080, 64'hf117b00000000000, 64'hc013839160acb56d, 64'h210420350df0a2d3, 64'hd13aa5d105cb56f4, 64'h18100e0739},{64'h3000240000, 64'h3099ca2000000008, 64'hbf8b6b015c5c8879, 64'h9e667e177ac005f2, 64'hc40209e38a011774, 64'h17d2ff70f7},{64'h200000014640800, 64'hf116bd8000000018, 64'h218e362c545ca90a, 64'hae5f37737ce1794e, 64'h4c48459152165840, 64'hb2c87381d},{64'h1400000043980, 64'h30f6a6e000001000, 64'h5840862c672cb889, 64'h5b0c185649f93f, 64'hc0b094d107ccf988, 64'h83f305b0a},{64'h194010080, 64'h4000, 64'h43899c18dba97200, 64'h35deda882ef48527, 64'h144c34a67e439687, 64'he04c51e83},{64'h51000, 64'h5ab4b02000004004, 64'hb40f55e65c3898a9, 64'h8a6f8a754ddee8ac, 64'h8d682bc71400152b, 64'h18f50b9311},{64'h1000008050800, 64'h3117582000003000, 64'h13cc6de45c427859, 64'h6a07b5a9bd456e5d, 64'h21700080c32c8591, 64'h1534505c00},{64'h4014611000, 64'ha6d5800000000018, 64'hdf0f342e54a8ac89, 64'hc509f87b4542defc, 64'hc742a4d38aa14275, 64'h1bf9c0165c},{64'h8000000000c0, 64'h80, 64'h6a4c6bdc98dae800, 64'h8b07a22cb483d747, 64'h8519537532a0b48, 64'h13ec019467},{64'h400800000030142, 64'h7138d64000000000, 64'h1d306d14562ee079, 64'h3b2360ecbdf6c145, 64'h4c735df5cd218430, 64'h698003be3},{64'h1805004000080, 64'hb138ad0000000010, 64'hd0f24035c288d91, 64'h29f014181a06d4f9, 64'hc0180fe18d3e0634, 64'h8386e10d0},{64'h410c000142, 64'h9abc0000000000, 64'hdff36a1656509700, 64'h75a191ec2405505f, 64'h347c50d0ae9501a6, 64'h2ba592644},{64'h501061000000000, 64'h30a0502298000000, 64'ha6c97e11572cad59, 64'h9316ce91d6093126, 64'h664b6199b66244, 64'h997ac5380},{64'ha000803000000000, 64'h30ab800000000010, 64'h14158da4d0a49499, 64'h8e2684b8840002cb, 64'h2848e65a7239734, 64'h2893400f0},{64'h14040980, 64'h500000000000219c, 64'haac99ca8d63cf1b9, 64'h350a1706406d5a57, 64'hd41a8004eeca9678, 64'h16b56a91dc},{64'h10000000, 64'h11605c078000008, 64'hcb90be164c000000, 64'h5fcb88702f4f2, 64'hb8870e66c0dc9b90, 64'h1940305a79},{64'h100c04000000000, 64'hb09ac1e000000000, 64'ha44c6d268bd96203, 64'h4004890148a40488, 64'hed69e9c2cfa704d6, 64'h7132},{64'h609000000020000, 64'h2b612c7200005180, 64'hcad134da57d0d789, 64'h2e05ccb12278570a, 64'h5d20784c81b30124, 64'h14e4bbed0c},{64'h500800010660800, 64'hf000000000000000, 64'h1d175ceaab44b20b, 64'hcf9d6366d0c82, 64'h74174aa4432a99a0, 64'h86475668c},{64'h410000000010000, 64'h9bd82000000000, 64'h4b0a5c1a47800000, 64'h8510a19520e170ca, 64'hb453e21da61905dc, 64'hf88765a64},{64'h5000000000200c0, 64'h30bbb94000004080, 64'hdf937daa8044b249, 64'h30740090f43a43d, 64'h1042e7461600c010, 64'h386d1cbce},{64'ha000000000011800, 64'h3117ce1590002010, 64'h6e01761aa05c9859, 64'hbd1726f599f2da3a, 64'hb7d00b0160005c9, 64'h18151e6fb1},{64'h6010050000000c0, 64'h30e6b02000001100, 64'h1491bce06958c9b1, 64'hc438b31029318433, 64'hc45ced3173148394, 64'h17d6ffda6c},{64'h418020008000140, 64'hd5000000000000, 64'h358bae28fbc49300, 64'h736ad359262f601b, 64'hd4624afe692a783a, 64'h6baf76609},{64'h8000040, 64'h9a800000000000, 64'h9f51a2ef342a0000, 64'hf75b12913e8a42c3, 64'hec0e81e03a078870, 64'h33a7b0ce9},{64'h300000008040800, 64'h2ef6b99598000000, 64'h8610881045248ba1, 64'h68142c336a3ac2, 64'h39a54fe5a0585028, 64'h8621957a5},{64'h10000000000c0, 64'h8000000000001008, 64'h178266d43d7672, 64'ha70b629c5905b0c7, 64'h402d8a75f91c0380, 64'h1bec7054d1},{64'h20000500c000000, 64'h1402c2000001010, 64'h1fd16ce4cabd3000, 64'hb2ad5715be07f4f8, 64'h417063546a0017bc, 64'h2877d5439},{64'h1010000000, 64'h17aa69308002014, 64'hb596261a57017800, 64'he34ef5a56b1e3368, 64'h28b21c250b28ce2d, 64'h1bfc8a0ff2},{64'h101003014060000, 64'h6f58bc2000000000, 64'h13601b6124cba1, 64'h5809b16044c862cc, 64'h4c51e8e06b4e0544, 64'h14996551ca},{64'h410000000010000, 64'h1750000000003000, 64'h74897da249a88d41, 64'h30606001c0506654, 64'hd42c5dfba6654434, 64'h8e72b2000},{64'h508004000000080, 64'h110ac4000000000, 64'h8577bad24d54000, 64'h3619acd866b05069, 64'hbc1cc3099a000117, 64'h1110b2183},{64'h200460014000000, 64'h5000000000004000, 64'h2791ace4ea256ab9, 64'hb704327802ad516c, 64'h5086c000af4376a2, 64'h74b74b52},{64'h1404000011006, 64'hb0582908000000, 64'he9308d685c4c9700, 64'h911c5dc5b7ac927, 64'h4ce99770094244f5, 64'he01600a27},{64'h101002000000000, 64'hf0c43212865180, 64'hdfcd4cd686000000, 64'hb5269d71680530a6, 64'h84ecc0b32d4474, 64'h43c5196a0},{64'h40, 64'h16a800000000000, 64'hd8179e1ea8d1a000, 64'h981309c197000675, 64'h800781301e04d950, 64'h1f8a007e2},{64'h518000000000000, 64'hf0f6b98b4a902010, 64'he2d48062590ef814, 64'h153812c87691480, 64'h304c789c808610ca, 64'h13d44c18b1},{64'h404000000144, 64'hb160482300000000, 64'ha4699adf185c98ab, 64'h42481109b402e0ad, 64'h1d6040539eb1c54, 64'h1963180841},{64'h418000008000040, 64'h1ed5d44000000000, 64'h7d154d090069861, 64'h3605d2784f09270b, 64'hb8046d193c4d80f9, 64'h100931264},{64'h400000000000, 64'h1000000000000000, 64'h22cf5c53554dd4bc, 64'h150000010c20410a, 64'hccecaf31550559a4, 64'h460003b2b},{64'h10450000, 64'h5b17d8400000000c, 64'hed4a86e44288c59, 64'hf21172161ec000cb, 64'h98932231a688c699, 64'h1bf83c0ed4},{64'h100003010000000, 64'h5824000000000014, 64'h2e4d8bdc585c8959, 64'h70077704e11a5667, 64'hb93ae340dc9d5c26, 64'h13a8001a71},{64'h301400000200000, 64'h3170800000004100, 64'h88be75a2c8e69, 64'h37b2e66221b256, 64'h848f6211f1b64b88, 64'h3751ec5c8},{64'h8053040, 64'hb141000000000010, 64'hc4d0b61756bcb851, 64'hed18997c2447b8a5, 64'h5d98e9c4e8cc14e2, 64'h2653},{64'h0, 64'h30b0800000001010, 64'ha64e981f71349089, 64'ha21c028322990cc, 64'h94338651f019d4c8, 64'h6be7b5391},{64'h40000000000000c0, 64'hb138bc2c08000004, 64'h149585d746c9c04d, 64'h135a024d9733b4fb, 64'hef3101350e24d9d8, 64'h1650530cf9},{64'h4280060080, 64'h2b16cde9b8000080, 64'h16d240e86c399881, 64'h778e02ed954a72c3, 64'h5d0001760041ae, 64'h10cd0c8620},{64'h5100010000, 64'h1215c3500004000, 64'h94f5e1cc9a89800, 64'h7094f0a82dc4708e, 64'h2922922244001b94, 64'h1842648a9},{64'h400018000104, 64'h5c9bdaa000000014, 64'ha22a23164c4cd869, 64'h310490e4db039489, 64'hf64503946b7089c2, 64'hb286b1779},{64'hc0, 64'h2c1000000000008, 64'h91d14e110c4db57d, 64'h48514120b4e8a5ad, 64'h383aa472cc1d53b8, 64'h1155},{64'h200000004000140, 64'h6f3880000000400c, 64'h4192855cb0308f69, 64'hb1b60dd84d483, 64'h3147502608030268, 64'h3add35270},{64'h1400000000000, 64'hb1583d6000001010, 64'h5a576893404cb80b, 64'he95d27918316919a, 64'hec110005a7791832, 64'h195c3b25b0},{64'h4014060800, 64'h3137deb60b063008, 64'hc2c932c10c44d205, 64'h91005cda1d4cde66, 64'h716e2b6722cd001f, 64'h116ff219b},{64'h501000000000080, 64'h2200000000001000, 64'h584b6b2d77a4b871, 64'h332660d16aed813d, 64'hb17d6d80170d0b09, 64'h36be2b24},{64'h408000000000000, 64'h137800000000000, 64'ha115ca0abb53500, 64'h2ef2d4858284f8, 64'h169dd3dee0a13b8, 64'h8627d5ee4},{64'h1000000000, 64'h1d30800000004008, 64'h157ded04d16851, 64'h7d03a1604c01d0b0, 64'h1c0d802fa0005ad, 64'h17bf2f5a36},{64'h10a0004661000, 64'h169a41408000000, 64'h59522d5c68accd00, 64'h491319ea52789e5d, 64'h5c260df03d077252, 64'hb394a47e4},{64'h1000000000, 64'hc0000000002180, 64'hb4b6e22a85d2800, 64'h7c5a65a82102d2f6, 64'h616b2e00b00010cd, 64'h1c66928991},{64'hc00000240080, 64'h30e5deb400000014, 64'hdf922b2c48b4b899, 64'hf1085cb25951270d, 64'h8049a1f75987c8a0, 64'h4f8000a10},{64'h18020100, 64'hb1a04c08005184, 64'h86158c2e5c348f00, 64'ha838b8144f58f0ff, 64'h30000003206289b4, 64'h1bec209272},{64'h219400000040000, 64'hb0800000001000, 64'h157baf3044b800, 64'hd01a6b50f1ed500e, 64'h24ecef3947b40f9a, 64'h466bd5700},{64'h300001000040000, 64'h3120800000002000, 64'hb54bb61e98cd5504, 64'h3468c4d04361b45c, 64'hf493747447b5469d, 64'h1e62f264a},{64'h44180010000, 64'h5a00000000000014, 64'h1e4f5de2a9daa991, 64'h348f2cb0e140054e, 64'h3d67b044eb1ba186, 64'h3d32b06bb},{64'h118000000000000, 64'h8, 64'h96cef242ecc00, 64'h602e3c9560986322, 64'h910e2ee62a713a2, 64'h1611935bfb},{64'h30140, 64'hc227800000006010, 64'h8056aa5145c22074, 64'he643a00176d0e16d, 64'h50f30000ca7550e9, 64'h5be9a1297},{64'h101005018600000, 64'h9f1638290000001c, 64'hcb90bcaa4154b859, 64'h11d9ef68186533, 64'h3032f3b2136f884c, 64'h180000a3b},{64'h100, 64'h1b800000000008, 64'hba4fae28b0350300, 64'h3f002bdd7b8000a7, 64'hec0003c07e0045d8, 64'h17503c5132},{64'he0010a0100000000, 64'hd0d4d26000000018, 64'h78d0585c78bd92b9, 64'h31e5678d96314522, 64'hfe4280002703e00c, 64'hf21d61410},{64'h8c00014061100, 64'h3000000000000000, 64'h6e09662f344ab4b1, 64'h405391012042ac81, 64'ha522e4aa45000e10, 64'h1192e10daa},{64'h400001000051000, 64'h8000000000000000, 64'h44095e2171c49342, 64'h6609c00017439c80, 64'h802064548a138b3d, 64'h1239112b23},{64'h800000000000, 64'h127b9a000000000, 64'hd975a62a0a2c300, 64'hf40014547a02c, 64'h9ce90160eb1e80b0, 64'h1b8271280},{64'h4000000144, 64'h30b4a2e00000000c, 64'hb6327d58a0b490b1, 64'hbf60e2fc0000010b, 64'hfc1da660769980ac, 64'h83e6665b2},{64'h400000008010000, 64'he0300000000000, 64'h15915cda97864300, 64'h755d31519b45456c, 64'h5bfc570ae1d4610, 64'h8f0000773},{64'h402180000100, 64'h3159c5e000000000, 64'h2acdbb816c2c9041, 64'h91ac22c4960b1173, 64'h356e4ac6692c57ff, 64'hadb8d158e},{64'h41000, 64'h30b4800000000000, 64'hdb137d5576c90105, 64'h18267e00626d8a16, 64'h4c812f74040010ca, 64'h14b3e67cc},{64'h0, 64'h4800da000001010, 64'h753be12b545d0b3, 64'h365344b94d000051, 64'hec000000c2a693e9, 64'h13ee7e1af9},{64'h611401010000000, 64'h9370000000000000, 64'h119e24fa2cb883, 64'hc60153b40ec931a0, 64'h4433d808cf460bed, 64'h4a1c60283},{64'h4094000000, 64'h62bb000000006100, 64'h44f982a54289849, 64'h4a9275e42e839072, 64'h482e1781462a809e, 64'h29d678b80},{64'h18001010061140, 64'hb0bbdaa000000000, 64'h124a2b1ae9d0b879, 64'h4a0e15dc53ee48b7, 64'h916b570aee590be4, 64'h1bf9cf39e6},{64'h800000000140, 64'h14000000004000, 64'h4b8e7cd2b55cb100, 64'h674204d89b06708f, 64'hd09793443f4c08a4, 64'h1361925e4},{64'h400002000000000, 64'h8358800000000000, 64'h1b537d1776aaec4c, 64'he55aa228c406d592, 64'h4544832122854e, 64'h251893120},{64'h1010000000, 64'h3137dea00000000c, 64'h9a2a56121b889, 64'hd5091bf16b2fc008, 64'h2004d2d25abf1686, 64'h9680544fb},{64'h301400004040000, 64'h309b000000002000, 64'h137d5a874560a1, 64'h269aa026c2b630, 64'hb1a3c2a019000000, 64'h117e360f4c},{64'h71000001000014c, 64'h30a0800000001000, 64'h336bb01a7a8a7849, 64'h2c3c99d0c38002d3, 64'h88116cfcc2188313, 64'h3d5886501},{64'h3000000000, 64'hb09a000000000004, 64'h11561eb84dc21a, 64'h32000000e983410a, 64'h311080c40488598f, 64'hc9c355850},{64'h10000040, 64'h30d5bd8208000000, 64'hdfc0762961d48989, 64'h5c0698763c00021d, 64'he56789b136001543, 64'h4d8797021},{64'h10001000, 64'h200000000000000, 64'he289a2ef15350e64, 64'h16b000df73bbde, 64'h2ea8e43c0010e0, 64'h2f38b5260},{64'h1000460100, 64'h309b800000005180, 64'h2150b39844349851, 64'h7e1770064c6d80b1, 64'hb4f22c25b0b041fd, 64'h197eead844},{64'h400c00000020000, 64'hd5302000001000, 64'h115e1cfa82f800, 64'hfa0608a996440000, 64'hc266e25250c55b9, 64'hf24433ad1},{64'h301000004460140, 64'h5f51000000000000, 64'h38138e1265b60091, 64'h3851022140005b, 64'h11949c0b1270000, 64'h4e0011c20},{64'h600000000000044, 64'hb000000000005010, 64'h91f55a5a8782f802, 64'h3cc2ecf30bb2cd, 64'ha849dd96d4799b50, 64'h4fd11841d},{64'h402000000000, 64'h159800000003010, 64'h61d27d1cb8349800, 64'h662cc1c03d4bf2cc, 64'hd89318f3a763c0b6, 64'hbd5b1191},{64'h440010000000, 64'h3110d40000000000, 64'hb9e1b77c93661, 64'h651a72fe3d03d6c0, 64'he01f2784cdcea2bb, 64'h3da4b07c9},{64'h62000000000, 64'h8a400000000004, 64'h1c11b61696aaac00, 64'h696d21c0b0800162, 64'h75b48200af47a617, 64'h388205bd5},{64'h100000000001800, 64'hd4d80000000000, 64'h179a22c9516200, 64'h2a2c417c58d348be, 64'h705661d548874b11, 64'h100860548a},{64'h4100000000, 64'hdc00000000003004, 64'ha6969a6119350f52, 64'h19bd6e3cf4b8f701, 64'h95532da0000014e6, 64'h865ea67da},{64'h201404000010000, 64'h1359dc2000006180, 64'hb331a6c4898a1, 64'h200401314d44c126, 64'h813ec4c0cbcd0f34, 64'h14d67ea6f0},{64'h3008000000, 64'h1b000000000010, 64'h79136d62b93c9800, 64'he4029864f22145f0, 64'he57ca19235170e35, 64'hbc09f65fb},{64'h40000000c050080, 64'h42f0000000000000, 64'h5a4dace91baecc42, 64'h1c1554717bda40bb, 64'h1e45ca12000bb9, 64'h10d1e24340},{64'h2000000000, 64'h7000000000000004, 64'hb4c84aa2e9c2e00d, 64'h1200000032aa60ca, 64'h6456000158194256, 64'h98ad439f8},{64'h110000000000000, 64'h30e6000000000000, 64'h17aa68fb2e2302, 64'h794bc0009b44e000, 64'he89a52fb12b316fa, 64'h27ae00929},{64'h14000100110c0, 64'h92e0000000000000, 64'hbf1192c2fc548882, 64'h9d4b56ac4adcb, 64'h21a412f48bcbc978, 64'h199000313d},{64'h460000000080, 64'h106cc3700005010, 64'hc8cf2a1646000000, 64'h5d271d7e5965ab, 64'hd99613725bb5ee38, 64'h1bd2b04f4},{64'h519040000010000, 64'h3000000000000000, 64'h10acd696b2e091, 64'h1f50c96c15c62100, 64'h401de36877b47432, 64'h2aa900aaa},{64'h6000005080040000, 64'h1750800000000008, 64'h4191b62139208a49, 64'h62bd60002a5eb068, 64'hca451072047983ac, 64'h196dd44ebc},{64'h6000000000000000, 64'h2b000000000010, 64'h32527d6ee6a58100, 64'h9b000000b10c92c4, 64'hce3cafe2563250f4, 64'h17bba871bc},{64'h20014400000000c0, 64'h7111300000004000, 64'h80957de8eb351849, 64'hcc5b83310eadc5a1, 64'h75d8cc5ef26fc38, 64'h14f850f3e},{64'h2000000100, 64'h200000000000100c, 64'h36516ce4cad2e049, 64'hd15b00013a0d103b, 64'hd5698d11b49b1474, 64'h2f4d25299},{64'h4000000000000000, 64'h1c9a800000000010, 64'h7fd47ae4c0b491b9, 64'h29036000bf62a454, 64'h6221812052000090, 64'h148001a37},{64'h2200c00000000140, 64'h30c0800000000010, 64'h2d95bd9c88b49091, 64'h459891121fe073, 64'hf724b70632dc4e0, 64'h710000251},{64'h4000400000000000, 64'h100800000000010, 64'h13ad1b77890300, 64'hed6d425dc1b6d706, 64'h473d9d71394608c0, 64'hde76ff4},{64'h801000040000, 64'h3120a40000000000, 64'he34d9e295b3e3061, 64'hd03ac00033de6da0, 64'h20372343b38d1b56, 64'h1c70000dcb},{64'h400010600144, 64'h308b800000000000, 64'h59b15d945634af91, 64'h8011549b258320db, 64'hb03b79f31f0f9c0b, 64'h1983273ed},{64'h110000000000000, 64'h1af1000000004000, 64'h115c2a94069851, 64'h886cd001b487c01a, 64'hf13c43eb1ee10c81, 64'h2f820e21},{64'h4000080, 64'h140a80000000010, 64'h1809b3dd182c9500, 64'h3f6d30003003f2c3, 64'h80c7ae25c4adc300, 64'h38d2b0f51},{64'h860004000000, 64'h3158ac0000004000, 64'h1485daf7053861, 64'h712c546c8e1662cc, 64'h75c407143ba92630, 64'hc4460f105},{64'h401420000000080, 64'h116800000006180, 64'h1313852abb288c00, 64'h2337c000100243d7, 64'h94066a6c43b6adf0, 64'h87deab0e0},{64'h4400000, 64'h140dc0000000000, 64'h158ae0a9000000, 64'h8a041cd2264a766e, 64'hb5c5bad5f25e1c5b, 64'h19c3123cae},{64'h200000000000040, 64'h1ae1282000004000, 64'hb5164a1f51b23059, 64'hb8433001492d43c9, 64'h9d7ce915b4000f12, 64'h1c5f80702d},{64'h4280000044000c0, 64'h680000000000e000, 64'h33558dd2b5021869, 64'h922395de848003a1, 64'h31615e4b24431539, 64'h1d84664356},{64'h800000040046, 64'h90800000000000, 64'h4db4bbdcb8821800, 64'h1496138206df0cb, 64'h13c24e4338750f2, 64'h16a67f4fe0},{64'h400000000000, 64'hc600000000002000, 64'he3896a9f183240ac, 64'h262000b0b8e26c, 64'h88ae8005ad488910, 64'h27cbc1785},{64'h100000000040000, 64'h217a800000000000, 64'h1462ed2c248a79, 64'h5df25256, 64'h5a4536658000cb8, 64'h1994011840},{64'h300004000050000, 64'h70b4800000000000, 64'h18db05d51021851, 64'h38f0005fc570ae, 64'h17565c0f8155334, 64'hf80074460},{64'h6000005004000000, 64'h309bbc4000004008, 64'h75152d82dc389852, 64'he650d8510fc98208, 64'h430cad3432b982be, 64'h3dd070aba},{64'h400000000000140, 64'h4400000000000000, 64'h624f6c593726c1bd, 64'h7f126000f5e7c163, 64'hfc105920fe255330, 64'h6527d3241},{64'h8000002, 64'h128000000000000c, 64'h58af961cb8aaedac, 64'h8a5fd0340698a193, 64'hf0b9b342e65219a1, 64'h15e31e751a},{64'h803000040940, 64'hf158d26000000000, 64'h9d0d4c18f705180a, 64'hd819961dc7edcd35, 64'h1372c243d74dc3e, 64'hc99923a67},{64'hc02000000000, 64'h4200000000004000, 64'h174a5bd3345d808b, 64'h38052a2c00000518, 64'hb69471b5ce068f, 64'h4a7172da0},{64'h1001100000006, 64'h3120800000000000, 64'h6ef4c54d64c96b9, 64'h12bc65b52e16d455, 64'haca60000b97fc14c, 64'h13c9eb4f27},{64'h400000001000, 64'hf000000000000000, 64'h8753655325a28a03, 64'h40a7a512514af0, 64'h404c01016f878000, 64'hf60003d80},{64'h1002180000040, 64'h30d5800000000000, 64'hb6889aaf27d89803, 64'h7bac82d16d068707, 64'ha4b383915975e8c6, 64'h1550690d2b},{64'h101040000000006, 64'h2e00000000000000, 64'h75ab6e253626aaa2, 64'h7005f834a035a1, 64'h94376253138d2000, 64'h1b686a0d48},{64'h300004014020180, 64'h7000000000001000, 64'h5acbab5345490099, 64'hb725b4e53d56b5f9, 64'h1cfd607062dc97c, 64'h19d3b6d60},{64'h1000020000, 64'h117800000000000, 64'h4acd9e2a9bb94000, 64'h8f2684b43e5332c4, 64'h320624c85, 64'h30ab80000},{64'h40000c040000, 64'h7080000000000000, 64'hc917bab395ae20a, 64'h3231f374315340c1, 64'h209a0bb5c5030978, 64'h198bb238e},{64'h200000000000040, 64'hf0d4800000004000, 64'h34d78a190aaa605b, 64'h5a048925248002cd, 64'h1c44d4500905402, 64'h1ac251a80},{64'h500004004000000, 64'h8000000000000000, 64'h2f137d1576ba304c, 64'ha337dc485e0a3162, 64'h3cc5371614c4dc, 64'h1c58532f20},{64'h300000000000000, 64'h558de8000000000, 64'hd4bd560827872, 64'h37c61db39be02a, 64'h49d6c6e1a436c370, 64'h19c4167003},{64'h2000030000, 64'h309b41a000004000, 64'h28d29d5540ac8e79, 64'h181460014958c5a9, 64'h8911a2243b10d5, 64'h694a41dc0},{64'h400001100000000, 64'h7000000000000000, 64'h2f51536f24b1ee0d, 64'hd6cf2330630bd198, 64'h21e4f219984c96, 64'h1278c718e0},{64'h4080000000, 64'h717ada6000003000, 64'h7b49a2a4f1011803, 64'h1ebca000af9eb2c2, 64'h702e004e6, 64'h1705ee4ff0},{64'h3010000000, 64'h1c00000000005088, 64'h79d7926d4054b879, 64'h2c6d571ccb80064e, 64'hb9c71ee71c000917, 64'hf3d379797},{64'h18000000020000, 64'h3000000000004000, 64'hcc4bbb6360b08e9d, 64'hdb07cc1ce3c3e1a2, 64'hc09bcc2c8e36d238, 64'h1c7458484c},{64'h102000c000000, 64'h2a90000000000008, 64'h720b9ddf68b95091, 64'h44fb98240000af, 64'h1c3b00007da23728, 64'he49a30fb4},{64'h460000040000, 64'h25800000000014, 64'ha2d0a4ee9430b800, 64'ha0fe18db4c7c0c4, 64'hf486079433757735, 64'h7107c0e39},{64'h200001000040000, 64'h7120ac6000003014, 64'h27896d628658b3b9, 64'h370e20001fc9e0e2, 64'h5ac96376688c83fe, 64'h13ef2f0c12},{64'h404000000080, 64'h317a800000003000, 64'hb60e48244b349179, 64'hd238a3646c0005b9, 64'he984d2e79c038c, 64'h16f67509a0},{64'h41940, 64'h5b71800000001000, 64'h51d48cd2f1324051, 64'h106d8899, 64'hc9049314124000, 64'hc9c4946c0},{64'h6101000000000080, 64'h7000000000000014, 64'h118d4bd8ec06f851, 64'h46432000f1846519, 64'h7ab6e175f38659c4, 64'ha69eb3cb1},{64'h400000000c000000, 64'h3000000000000004, 64'h44958dded901184d, 64'h44d840b6d1237a, 64'he6330000cc3c4de8, 64'h10f1b93d79},{64'h3000000000, 64'h1c00000000004100, 64'h78957de09b226161, 64'h16a000b22aa072, 64'hf034a1a4342f0ebc, 64'h33579bd92},{64'hc0, 64'hb0f5b04000000008, 64'hdb4dbba9208eb805, 64'h408e41c03905b5, 64'h4574c6a000001020, 64'h88000d30},{64'h6000000000000100, 64'h2ab4342000000004, 64'h5840862971025899, 64'h9d80071d, 64'hff12c6e7521b9d48, 64'hb013c0d55},{64'h800000000040, 64'h20f6800000000010, 64'h441a62e80053871, 64'h5e7482f9d20002d7, 64'h7c0380070901cc80, 64'h600120031},{64'h1400004000000, 64'h289bc0000000410c, 64'h89e2255b08f91, 64'h30269cc06f0ae15c, 64'hcc8e3140ab64256b, 64'h3d63dc90},{64'hc00000010000, 64'hb0000000000000, 64'hb5516ceb0b328200, 64'h9a566482, 64'h9c1295d711a9c6a0, 64'h19ed44b65},{64'h100002000000000, 64'hb0c1c0200000400c, 64'he0556ad2fb82d812, 64'hc90a6e7524c00314, 64'h2c6a40d392001405, 64'h655a804b6},{64'h3004042880, 64'h7120000000000000, 64'hc20e4c6c45ddb899, 64'h2f3de8c540de73, 64'hc86933d0a7cf5c5c, 64'h1c093726e4},{64'hc000000, 64'h26000000000000, 64'h260dbbd2b5226100, 64'h1b70b0df42c052, 64'h5200031a000000, 64'h150ed1320},{64'h800010600000, 64'h2aabb02000001000, 64'he43762c44093899, 64'h5364b3c800500, 64'he88d43a2259b12f8, 64'h526814a00},{64'h200000000000000, 64'h8600000000000000, 64'hbbb6d04d1e112, 64'h7d020df52307f48c, 64'had3fde447e000083, 64'hb108018f7},{64'h400c00000000000, 64'h269a850000000000, 64'h19d47596d1409289, 64'h8e26819c9a24748e, 64'h94085eb703914f43, 64'hf74683d87},{64'h860004000000, 64'h3149444000000000, 64'h2c979a6afb356a04, 64'h316590012100007c, 64'hccf740071d72e693, 64'h1941ee3cc2},{64'h1100030000, 64'hbbd86000000000, 64'hb50956054c06188a, 64'h47b460001f4b716e, 64'h1d3d25d18e0006de, 64'h16b2b94f23},{64'h200004000000000, 64'h2ce5800000001000, 64'he4974a14d60658a9, 64'h835cd001c935a216, 64'h3bc00204e105bf, 64'he4c636d80},{64'h300000000000000, 64'h400000000004000, 64'h36d4ade2a7d9c149, 64'hd86683603e4db176, 64'h1464d11a23545d8, 64'h30cd10000},{64'h40000010c000040, 64'h2d20000000000000, 64'h34d57de299b52e81, 64'h37c6534c100000e3, 64'h845dcd909a0019a6, 64'h6c8211b20},{64'h300800000000000, 64'he1800000000004, 64'h9a2d576a26000, 64'h92000bf8002f4, 64'hf426cbd3a7328650, 64'hc00ca4eb2},{64'hc040142, 64'h3120000000000008, 64'h64af4c1656d088b1, 64'h46d1dc51d6d179, 64'h343c29b0938d10c8, 64'h23a9b2df5},{64'hc05000000004, 64'hd4860800004000, 64'h5b755e26563cb800, 64'h120000000000008d, 64'hc87906d3d71b4376, 64'hb46d43c3},{64'hc00000000002, 64'h3000000000000000, 64'h6f6d4bd511017803, 64'he200038899225, 64'hf8868be0cd1c48f8, 64'h4d00023e2},{64'h10006000000010a, 64'h1a8a800000002000, 64'h33327d185c28b059, 64'h2f662c09bd06c17b, 64'hb3fb1435ba702a, 64'h16df814620},{64'h30000, 64'h400000000000000, 64'h6f51aa9b39268104, 64'h660006f5c8400278, 64'h85d53a944b198dd8, 64'hb12a654ca},{64'h3000000000, 64'h9917850000000000, 64'h95aa70b82c26c, 64'h1a00eb6d6dab253a, 64'h79a129e43478dd4e, 64'hb672f684a},{64'h2000800000030000, 64'he321000000004000, 64'h2553ad1766a92c73, 64'h6b462001d2714384, 64'h7e4a89300f000e10, 64'h2c5b91811},{64'h400000000020040, 64'h7000000000000000, 64'h59928e18dbc13605, 64'h661b548e55f15d, 64'h83e4a48a8d4000, 64'h1650130260},{64'hc00010000000, 64'h30a4800000000014, 64'h953406f5035c279, 64'hff2a4d400d350, 64'h98000005050004f0, 64'hc5b824fb0},{64'h100, 64'h44bb850000003000, 64'ha6016c4e184d, 64'h20e0005f90713d, 64'h6009919e264e4c, 64'h1cf4996fa3},{64'h4000000000000100, 64'hb000000000000004, 64'h1cd4be4eaae8c12, 64'h781965e0658085b1, 64'h69600067b32c041, 64'h5592c26fe},{64'h200000000001800, 64'hc4800000001000, 64'h33d144e17ac9f400, 64'h47c000c942ccf2, 64'hd88a66e4c03701d0, 64'h156761b69},{64'hc0, 64'hb100000000001000, 64'h40992d577d9a20b, 64'h75546a70082a2505, 64'hcc1d4000209d5bea, 64'h140e734ea9},{64'h100000008600000, 64'hb1415c4000000000, 64'h9dca5c6b39292f83, 64'h22021df60000048d, 64'ha8f646815c2b13d1, 64'h5782a3d20},{64'h501060000000040, 64'h30b4b40000000008, 64'h918e7a06ac5cb089, 64'hce6a88790a09d48f, 64'he834e1e1797bbaa0, 64'h346403d95},{64'h5100000000000c0, 64'h4200000000000010, 64'hcb0bae1b49c232ba, 64'h383dd1dd8b800663, 64'he0354dcc768e9963, 64'h35b280232},{64'h101000000000086, 64'h30b1800000000000, 64'h2df1a6209bbd0e99, 64'h70606dad81b395, 64'h13d5ec0dd001ad8, 64'h16b76d3d80},{64'h20000500c000000, 64'h2ad5000000004000, 64'h2b9248410c029899, 64'hd10c7345b4800725, 64'h188678015ee04c84, 64'h94d615ce},{64'h800004000006, 64'h7131444000000010, 64'h2eeba61b47dd4e02, 64'h251b1094150001b7, 64'h5c088b21a30846c8, 64'h88b20673},{64'h408005000000000, 64'h30d4b10f00000000, 64'h635058825c4493a1, 64'h331940ccc9000324, 64'hcc12cd997a41c6a4, 64'h839050430},{64'h100000010000000, 64'h12038200000200c, 64'hb4484be2b9d2f600, 64'hd80a72e05c2d12da, 64'h445ec00170a68654, 64'hc054e2f73},{64'h101000000000000, 64'hf000000000000008, 64'h157de6ea59208a, 64'h9b4281b400000026, 64'hcc3c61e1a5700e18, 64'he181446b3},{64'h500000000000000, 64'h309b4c0000002010, 64'ha74f8a1b20896381, 64'h995a25b0b61430e2, 64'h8c526a30db2f968a, 64'h89c72133a},{64'h300002000000000, 64'h903c7600000004, 64'h9fd3ad21192eed00, 64'h45800038f2f454, 64'hc5f61f0000008fe, 64'h14025721fc},{64'h2180000000, 64'h3000000000004014, 64'h66574a2d19556169, 64'h2692a000de895208, 64'hc6861ce128739c0e, 64'h4050c2c58},{64'h300005008040000, 64'h1a000000000000, 64'hcc0dbbe4eaa6cc00, 64'h9e2dfba09a7305b6, 64'h55d56e7566001c76, 64'hb400054dc},{64'h110003000000140, 64'h3110800000000010, 64'h46155dc0eb34b341, 64'hbb384e216df8807d, 64'hb14f7429e00010d5, 64'h1ae9191671},{64'h1000000001840, 64'hf000000000000000, 64'h14d772668aca2202, 64'h9337a6ed18f3192b, 64'h502a00018f2544a8, 64'hb39be2c41},{64'h800000030000, 64'h8200000000000000, 64'ha6929a5f182eec42, 64'h11b5a95ab, 64'h15532a5495314628, 64'h11707b45e3},{64'h3010000000, 64'h4200000000002000, 64'h1d8dbb1eb8212a05, 64'h846697269a2d55aa, 64'h31c237f180001c17, 64'h5547526eb},{64'h20100000c010000, 64'h30e1000000000000, 64'hb4174e18d8d57655, 64'h70302083ece196, 64'h886040809b267588, 64'h662e25a2b},{64'h10020000, 64'h81584000000000, 64'h982ef554da100, 64'h935e265cd0000, 64'h6d8004e0001510, 64'h13d22d0000},{64'h418000014000000, 64'h3000000000006000, 64'hdc8709950a4b881, 64'h374332654283750a, 64'h854de82932945518, 64'h23c004eda},{64'h8000000000c0, 64'h137000000000000, 64'h2ed58de8fb416100, 64'h94176000e61c36fb, 64'h351cc4eb2693ac, 64'h13c0001340},{64'h100c000000, 64'h3179000000004000, 64'h33c8609447b634a9, 64'h1e24986483ad548e, 64'h593aacc13c9d4f76, 64'h4d4afa10b},{64'h8000000, 64'hb0f60ec000000000, 64'h8e956ae975466103, 64'h386a9cb14e8d362e, 64'hbd7546a8335953, 64'h14f0d40da0},{64'h1404000030000, 64'h848a26a000000000, 64'hd7ba700c6d8ba, 64'hc671d703bf836da, 64'hfd3b0002c5000335, 64'h861054ec8},{64'h10030000, 64'hc400000000001000, 64'h84c54b656c00c, 64'he00f3580de550fe, 64'h4028650ccdd9bb, 64'h1c9caf1000},{64'h400000000000, 64'hf024800000003000, 64'hf8c1b572acc1c, 64'hab0305e012800028, 64'h1c3c157030680d0, 64'h6e5790300},{64'h4100c0, 64'h2141000000000010, 64'hcfd38a6c46a89279, 64'h261b30966cc33055, 64'h1c1326067ac24c80, 64'h1408000274},{64'ha000000004000080, 64'h2350816000000010, 64'ha6886e1cfb8a1861, 64'h9f067d506c000325, 64'h2e000001a4720e41, 64'h5c8cf04d6},{64'h10000, 64'h8680800000002000, 64'h4d0f8c269c02f8a3, 64'h9c2580005c4005a3, 64'h1ca0002584d4e00, 64'hb7f677280},{64'h6400400000000000, 64'h1e00000000000008, 64'h738a4b21103892b9, 64'h4a3dc7a4e70492d8, 64'h129659e43d510f70, 64'h238002297},{64'h200004004000000, 64'hec00000000000000, 64'h2b554468dbc27203, 64'h1b5a395cb661e630, 64'h151e1c1060001d4, 64'h57000662a},{64'h4040146, 64'h708b800000000000, 64'h87ed755561026b89, 64'h4590000842c021, 64'hc83a756880013a8, 64'h140495218d},{64'h500000000010000, 64'h3106800000000010, 64'h57ca60829c2c8ea9, 64'h5c245c4ad172cc, 64'hb4344e339d59d708, 64'h16e2b4055a},{64'h300000008000002, 64'h5000000000000000, 64'hb6f6bbe0b94db50a, 64'h5d14843611f661, 64'h80b443f2e6280500, 64'ha483f2ea2},{64'h10086, 64'h26d4800000000010, 64'h8c6f5c1c850e98a9, 64'h7c3ea1f1c45bd385, 64'ha83d9f30a888c2a0, 64'h8ce2a1718},{64'h410001000000000, 64'h10102ae1000000c, 64'hcc0f6e22c9a64b00, 64'h7f18ac559892e0f6, 64'hb8f64548000004ad, 64'hbf12f2cf8},{64'h5090030000, 64'h709ac82000000000, 64'h179d1761209141, 64'hc59a3044e55672ce, 64'h855353702200068c, 64'h170aa9164b},{64'h429801000000080, 64'h3036800000000000, 64'h2084aeaab38b3a9, 64'h722e46f4619bb5ab, 64'hf85941184330dc25, 64'h3bed127c6},{64'h1400010020000, 64'h14dc4000000000, 64'hb393aae2a93cb400, 64'h85195d6c046a25aa, 64'h91121fb17bb594e3, 64'h1c38005c58},{64'h4000400000000000, 64'h600000000000000, 64'h3a16bbe3342dacac, 64'h53032d4c0c911222, 64'hb6000001b90600c3, 64'h1c09c4f58},{64'h14400002, 64'h2880000000004000, 64'ha1714ceb7b3c9091, 64'h5d0dba8fc4b8806f, 64'h4d0000ec000e63, 64'ha49a0ee0},{64'h1400000000180, 64'hb016000000004180, 64'hb5558d1c45412271, 64'h1b0345670d90e3, 64'h7d0b91717d8793d4, 64'h395c4a2e3},{64'hc00000000000, 64'h4, 64'h57ca5b653abd82bd, 64'h670001963182c2, 64'hece89622f5000000, 64'h370002118},{64'h100, 64'h61a000000000000, 64'hbd96bb655130985a, 64'hf14520017b88037b, 64'h57f0006a9bf9149, 64'h17c0815f02},{64'h100864000000000, 64'h1400000000000000, 64'h6f508c9977a6ab45, 64'hce6e750e11d4384, 64'hc93b493709e5b4f5, 64'hb913a61e5},{64'h200400000000000, 64'ha40000000000000c, 64'hde084ae6dad2f602, 64'h137140003c000706, 64'hc04078b50de119bc, 64'haa301b98},{64'h3008000000, 64'h4200000000000000, 64'h944d961345daef44, 64'h9e0312d589aa350a, 64'h5151800510d540d6, 64'hbcd9367cd},{64'h3000000000, 64'h224800000000000, 64'hb9bed77323555, 64'h805a27200000019a, 64'h80610806a8000134, 64'h14d0005036},{64'h10000000000c0, 64'h3116800000000000, 64'hd68eb06481017361, 64'h2c6ce001c90001b1, 64'hb521000181000e45, 64'h8fa4226a4},{64'h140, 64'h70c48a2000004080, 64'h740096297c296341, 64'h5cc12517800197, 64'hc5ca5ec39c669d80, 64'h665c3c621},{64'h8000046, 64'h7000000000000000, 64'h5b309ca8b539f713, 64'h3dd70d7f00039d, 64'h89402585febe4254, 64'h1590005c8b},{64'h10201800, 64'h3000000000000008, 64'h147b968509ac99, 64'h7f133cc70f41c800, 64'h505e00e6fe0004ab, 64'h5e0c35012},{64'h800000000100, 64'h3000000000003000, 64'h138e6c60b0a08c49, 64'h5204e177, 64'h9486564689928270, 64'h16ca52ce2},{64'h1000004020000, 64'h4000000000005180, 64'h1585d345bcb853, 64'h5c30008bca023e, 64'h8c6b8004eb2f06b8, 64'h1246dc9b2a},{64'h80, 64'h3150000000004284, 64'hc8d678d45c30b059, 64'h7c6629e08b8e3467, 64'h419891a0f69e8504, 64'h14f4d4aeb9},{64'h4000000, 64'hb000000000000008, 64'h18535be956b2f28b, 64'h170f900117289514, 64'h8c3186100000111e, 64'hbc8004551},{64'h1002000000000, 64'h300000000000000c, 64'h5b0b6b2b7b522141, 64'h138400198dbb054, 64'hece180015fc04bff, 64'hb69452fdb},{64'hc00008040040, 64'h3000000000000000, 64'h812ab1eb8dd28b1, 64'h2002330c12dbd2cf, 64'hd03b8202d12f83a8, 64'h1a0775c30},{64'h1400004040000, 64'hc40a800000000000, 64'h59d16dd306208b9b, 64'h2e5e1419cb23f6, 64'h5c6e00020f891ae0, 64'hb50001b83},{64'h2000000000000c0, 64'h200000000004000, 64'hdf17aa14b60acf9c, 64'h9c2e44f800000545, 64'h5127815ad000748, 64'h5cd122eae},{64'h2000030040, 64'h7000000000000000, 64'hbbb6535060904, 64'hb46a71e40cc00223, 64'h791808746021c0c6, 64'h16e0876feb},{64'h3000001000, 64'hb000000000000004, 64'hd4bd937222b02, 64'h701b22b5c4dccdf0, 64'h580b536a60003b5, 64'hb889b0efc},{64'h8000000, 64'h1900000000400c, 64'h119a1a972ecc00, 64'h43d1f08e11b0f6, 64'hf48bcee18e4688c0, 64'h575625ad1},{64'h864000010000, 64'h4800000000000, 64'h26506beaea4ecb00, 64'h33458bd99cdc3386, 64'hd84092c3a38ef3ad, 64'h1813014547},{64'h6000400000000000, 64'he4c1000000000008, 64'hba516e2b7b266852, 64'h4530fd9bb0f278, 64'he2000005fd0fc000, 64'h103b},{64'h40000000c010080, 64'h3000000000000000, 64'h1343ad016c3c93b9, 64'h5c66f134ea77a385, 64'he01fc795f0001c58, 64'h1c204e2e5b},{64'h301804000000000, 64'hb0e5820000005004, 64'h32979a515105b889, 64'h5463299e304678, 64'hd00ae560a9a182a4, 64'hdf4cb4614},{64'h140000c0, 64'h3029000000004000, 64'hbd79a695b3da159, 64'h18b5c4e41a067f, 64'hc4188006ab204000, 64'h97d631020},{64'h1060008000000, 64'h30f5000000001000, 64'hb68bbb124c0ab499, 64'h391d6daa6d3724, 64'h16b00026f30a000, 64'h1696ab0a20},{64'h860000000140, 64'h10, 64'h73974e2aa65a6100, 64'h3e67c000f719e011, 64'h5bd381126b47f53b, 64'h1733165a3e},{64'h0, 64'h3a000000000004, 64'h734c6e22995ea244, 64'hf75c2ab4e69955f8, 64'h17f8005fc0017fa, 64'h4630},{64'h200000000030000, 64'h8000000000004000, 64'h14addd184a6165, 64'h39e000e2dd712a, 64'hf1404006fe038e78, 64'h1c5a701e2},{64'h1000180000000, 64'h301b096000000000, 64'h23104c80ac39f8a9, 64'hc3b846ed2c08f11e, 64'hc52a80135a09bfc, 64'h2780009e7},{64'hc00008000000, 64'hc0a80800000004, 64'h2a129aeb7b368f00, 64'h1f49587c4008609d, 64'h88ef8002cf18c31a, 64'h548a614b1},{64'h462000000100, 64'he000000000000000, 64'hb88cae2349dd287a, 64'h702431f03dae2659, 64'h455d0001b3a8e6be, 64'h13d2d65acb},{64'h100000008000000, 64'h600000000000000, 64'h86d565d2b522209d, 64'hc663929ac80045c, 64'h648d42620e099251, 64'h13399218e},{64'h3000000040, 64'hc538000000000000, 64'h7089a2da87a9d1b5, 64'h1802a17d8c0515, 64'h31ca41802a4bcc, 64'h3800},{64'h10000000c0, 64'h8000000000002000, 64'h8bd36be4ea8698ba, 64'h75040cc4df325057, 64'h1a04a66212980c, 64'hb6c494620},{64'h4100000000030000, 64'h30c1024000000010, 64'hd4bef153ab3a1, 64'hfc00000061f85000, 64'hd23bf6843e8cd121, 64'h11a0003270},{64'h100804000000000, 64'h1000000000000000, 64'h28c2ad1b89879, 64'h45484001229d9000, 64'ha86e400449908406, 64'hb54002243},{64'h400000014000000, 64'h7000000000002184, 64'ha2425a9e494494a9, 64'hd825921c31219514, 64'h1d21781c3285c439, 64'h89756aeb2},{64'h200000000c0, 64'h130400000000008, 64'h18515e1cfade9600, 64'h2e000047086713, 64'hbc3189010f8c2a28, 64'h5716d5bd5},{64'h200400000000000, 64'h0, 64'h5e94ab597c260b92, 64'h65a28c3e1691c2, 64'hd980d176a7471968, 64'hb517b20ab},{64'h0, 64'h808a8a8000000000, 64'h179a60b93d416d, 64'h882664b000000000, 64'h1808005f2d4c4d8, 64'h1ab08f11e0},{64'hc000040, 64'hc000000000002000, 64'h2a498a9f0431d894, 64'h3f4598a50122c387, 64'h21159f4456000550, 64'h18144a0941},{64'h4040000, 64'h202880000000000c, 64'hd7536d5947256ab9, 64'h992ebe6450737810, 64'h1027009012a15443, 64'h1bea505d5e},{64'h200c000000, 64'h2c0000000000000, 64'h70d1bcde9836ce5a, 64'h9a0b9c1d9b9c5672, 64'h1880002f4001184, 64'h2749f1960},{64'h860000000040, 64'hf0a0000000000000, 64'h5cce4e2f1ad1960c, 64'h603ae264b9800679, 64'h30a59d85114d2180, 64'h65e8c2c8a},{64'hc00000020000, 64'h3015000000000000, 64'h129b68cba62b04, 64'h30000000e4400556, 64'h18dd12ed8c1ae2, 64'h1c9adb0f40},{64'h100000000000000, 64'h3000000000000010, 64'h1c8f54510126c069, 64'h550000e4072394, 64'h996b5a1228000390, 64'h888e137db},{64'h4000080, 64'h8600000000000000, 64'ha3084bab0bd1b65c, 64'h5e67d14c9e2263a1, 64'hc9459754467cdd3e, 64'h14380050e5},{64'hc01000000000, 64'h5400000000000008, 64'h170e7d5746b27744, 64'h7a2f4000d485c39b, 64'h3c4f8565ffe057fd, 64'h868cc5c94},{64'h4000c0, 64'h3017800000000000, 64'h156dd095c59205, 64'h39fdfee12ab3af, 64'h6e2e4000000468, 64'hdf0005c20},{64'h800000040040, 64'h0, 64'hc10aab584c0618a2, 64'h114c0046cf3c11f, 64'h505000b78, 64'h1a00000020},{64'h400003004000000, 64'h3000000000002000, 64'h2055ba22a98a5881, 64'h3343f9e83e3526a4, 64'hccb15e080000031e, 64'h54e734f49},{64'h400000000000000, 64'h303a000000000004, 64'h734a5ceb7b292289, 64'h9804cd70000005c5, 64'h40d0c442424131, 64'h1179d15ad0},{64'h400000000000, 64'hf120c02000000000, 64'h178a50e1b5e204, 64'h7f38e65ce1000180, 64'hf80000004dbf1c0b, 64'he580f7336},{64'h1000014410000, 64'hc760800000000000, 64'hc9d14c253409f8a2, 64'hc7717c06604c437e, 64'h69b10c85f12a7988, 64'h1cd00054ce},{64'h40000, 64'h303b000000000004, 64'hda11ab50c5c2e251, 64'h43e00151c0070a, 64'hb100009559d198, 64'hb38004630},{64'h1000000000000, 64'h600000000000000, 64'hb38863ed70c88281, 64'h424601fc638005a0, 64'h19689d6103759126, 64'h630004622},{64'h200c0, 64'hd418800000000000, 64'h14461ab7daec94, 64'h8a0920bd22c003b3, 64'h139b41094d090d2, 64'h2250},{64'h900, 64'h400000000000000, 64'hb88d9bdd2c40988b, 64'hfe1d4898ec619bdd, 64'h8a0005febe1122, 64'hfeabd2240},{64'h0, 64'h2600000000001188, 64'h174e22f72a4c82, 64'h9000000ea00023e, 64'h484a40000008e1, 64'h32571adf0},{64'h428c00004000000, 64'h7000000000000000, 64'h1426211101b8b1, 64'heb65b00000000000, 64'h4b4bca35000bea, 64'hbdeeb1120},{64'h400000000000086, 64'hb000000000006094, 64'h4ce056204c24b149, 64'hba65abd996a19603, 64'h3e52cc11820010c8, 64'h27f5689f2},{64'h403000000000, 64'h158000000000008, 64'hd8ba53a000000, 64'h8666cc191665b000, 64'hfdc211a457468556, 64'h8033a095d},{64'h800000000000, 64'h4200000000000000, 64'h129a5a87b1638d, 64'h6373319cbd862162, 64'h13b27b0139ece28, 64'h320000000},{64'hc00010000080, 64'h8018000000000000, 64'h8a8d9be3543098a5, 64'h82495800eba2c673, 64'h3c000006810004d2, 64'ha70004fe9},{64'h30040, 64'h8, 64'ha5c6f3a8518a4, 64'h6372600018f932e7, 64'h44108000000016f3, 64'h1082c519b},{64'h408000000000146, 64'h7000000000000000, 64'h74728d60b120ac49, 64'h90ea1b41802e041, 64'h401a796862025184, 64'h398cf0ee4},{64'hc000044, 64'h117a02000000000, 64'h72ab4e29574a6a00, 64'h235cd000000000e5, 64'hfa2612295cd45a, 64'h2c0002920},{64'h0, 64'h700000000000000c, 64'h1590409ea0c5801b, 64'h3be7784800021c, 64'h1000000122000000, 64'h50f2},{64'h5010430000, 64'h701b000000000000, 64'h7080be28474d72a1, 64'h10f5eae843f0b9, 64'he1750001b8b8843c, 64'he02ea11ca},{64'h0, 64'hc017000000002000, 64'h9ab04ac5d037a, 64'h775cc00000800000, 64'h53ae6000001181, 64'h486cf0000},{64'h40000000040000c0, 64'h3140800000004014, 64'he00d4ca05c099889, 64'h43003d0dc036d2df, 64'ha73d02e4ea0013ab, 64'hb57408fb2},{64'hc000040, 64'h0, 64'h69116ce95bb1c264, 64'h467759771d66a5, 64'h101f800218000450, 64'h17780039e1},{64'hc00010000000, 64'h3027000000000004, 64'hd493855570518859, 64'h7fd58e38005ac, 64'h400000739208cc0, 64'h1be9c345fe},{64'h400000000020000, 64'h3034800000000000, 64'h38577ce900ad00b1, 64'hd718e31580c98678, 64'h60276a6228001839, 64'h1a00002227},{64'h2000000008000000, 64'hc036800000000010, 64'hc11aad5775a0894, 64'h41663de80000070c, 64'h6ab3a212ee110220, 64'h1882f197e},{64'h4000000000, 64'h300609a000003000, 64'hbf0f8c2e945a6171, 64'h573200043301602, 64'h14000006bc010b24, 64'h11a6d17380},{64'h400000000000, 64'h302480000000000c, 64'h4ecb7c64e556f60d, 64'h30436e50243942d6, 64'h28b78003add04644, 64'h1b60004631},{64'hc0, 64'h4029000000000000, 64'hb9d3456d762e817c, 64'h642d20d41aae7515, 64'h14600006a11d7f9, 64'h308005180},{64'h20040000c000000, 64'h7100800000000000, 64'haa957de6ea290c94, 64'h6444d470000005b4, 64'h9c8a6de5ff09c139, 64'h17250f04e5},{64'h10000000040000, 64'h420000000000000c, 64'h878b8e1ea85aed9a, 64'h5149ddc0c89514, 64'head7bc3c85d978, 64'h1990382410},{64'h2004000000, 64'h700000000000000c, 64'h11104a1cfbca7605, 64'hc22fb5e80000013e, 64'hec47d7b0860ed75c, 64'h608b95d72},{64'h10000, 64'hf000000000000000, 64'he7dd098cecd02, 64'h750cb9d96f36000, 64'h8e8b6183971c23, 64'h2380023a0},{64'h440000000100, 64'h4101000000000000, 64'ha6b268c49e3ac, 64'hc6d15a50c60f9, 64'h2000000235e13a50, 64'h158c804c3},{64'h65010020000, 64'h7019000000000000, 64'h9f89aae0aa4d5841, 64'h2a04dcc53be7e662, 64'h9d3fb964f75f2137, 64'h12824b728d},{64'h300000000010100, 64'h2000, 64'he4d54dd4b6ce3662, 64'h5d000116677181, 64'h4cec40038a9dc1d0, 64'hbaee76c87},{64'h410c00004000000, 64'h3157800000000000, 64'h3149849c4c015759, 64'h545bd451c9cc718e, 64'h68e042185941c2e0, 64'h2f33f67ec},{64'h400000000000, 64'hf000000000000008, 64'h56895aa11456f69b, 64'h8670c00000000229, 64'hd576800063a30333, 64'h1b58000ef5},{64'h300000010020000, 64'h3000000000000000, 64'h11449f002ee161, 64'h4858b11362c000, 64'h7d444864240002b8, 64'h488001187},{64'hc0, 64'h4400000000000000, 64'hb25375410c21415b, 64'h11c1642c800121, 64'hdc3b8005d21641d0, 64'h2edc35c81},{64'h0, 64'h30c5892000000004, 64'hdc937d032c2ae374, 64'h2ee891133723fc, 64'hc9754005ccb4db90, 64'h11906d1218},{64'h200000000000000, 64'hc039000000001000, 64'h1585d095ced473, 64'h658ca817000000, 64'h54f8670c0013b8, 64'h118f2d6d40},{64'h800000000040, 64'h3000000000000000, 64'h740d53a5348a0305, 64'h4e6876d853800701, 64'h84548214f5000548, 64'h116ad75ae0},{64'h300000000040000, 64'h30d5800000002000, 64'h30098a99485e6141, 64'h1e23c0010cdd6b90, 64'h1422400184324839, 64'h177d073464},{64'h2000000000, 64'h8200000000003000, 64'h117c92b83af8b2, 64'hec6ad10c21800626, 64'hf4e9912000001c0c, 64'h16cc0067c0},{64'h300000000040000, 64'h4200000000000000, 64'hde135d184c2ac26c, 64'h708000e2c68700, 64'h8647526a4001c08, 64'h1c100e3b11},{64'hc0, 64'hf000000000001100, 64'hdab90995af002, 64'h3c678c0db11d62ef, 64'h2d3e8684f6000227, 64'h18f87f342},{64'h80, 64'hc600000000000000, 64'hd0519c9cd62a81aa, 64'h4a70ad709e36c603, 64'h60800002c, 64'hb600070e0},{64'h4000000000, 64'h7028800000005000, 64'h129aaee1a28105, 64'h3273a001ca56901a, 64'h5412614641c404e, 64'h39c3673ca},{64'h200000000010000, 64'h3aa42000000000, 64'hb6b256539f100, 64'h7723809c1aeab5cf, 64'h14656700a1dc028, 64'h16d8050d80},{64'h1000030000, 64'h313081a000000010, 64'hf545c9822a291, 64'h1e0000008e61975e, 64'h21a18006860b413e, 64'h21f4},{64'hc04000000080, 64'h3000000000000000, 64'hc7b964c46a1b1, 64'ha20000005d83f515, 64'h80000011fe886e7, 64'h1994020880},{64'h200001180040000, 64'h2200000000000000, 64'h2d83a61550248b79, 64'hc185e00000c3166e, 64'h48bdc00510000614, 64'h188004dcc},{64'h0, 64'hf000000000001000, 64'h8955ca1596305, 64'h1aa28a514, 64'h8ec0018e468810, 64'h1744004fa0},{64'h6000004000010080, 64'h3000000000000000, 64'hcb1555a84c01d87c, 64'h204b4001a573168b, 64'hae62000500480865, 64'h1ab0001910},{64'h408000000000000, 64'h3000000000000000, 64'hc60f645d21d6e241, 64'h526a4cf9b20694fd, 64'he1f96800000e2b, 64'h1693946800},{64'h1000000600080, 64'h1218000000000000, 64'h4513baa359209815, 64'h5c5d174e00000727, 64'h1ce00054dd54863, 64'h1178007320},{64'h1005000000080, 64'h600000000001000, 64'ha8b105c3c98bc, 64'hde5d0481b692018f, 64'h14218002cfb9d10e, 64'h2f40067f3},{64'h410c00000000040, 64'h3000000000000000, 64'h8b935d5ec9029889, 64'h70d87800000519, 64'h1d68d75ddb77c000, 64'h4422},{64'h800000000000, 64'hc600000000004004, 64'h164a262e4c4c987a, 64'h4c0011642b602, 64'ha8450a512323c550, 64'h10e42b0bb2},{64'h200c04000000000, 64'h370000000000000, 64'h11c99556d858987b, 64'hff0da0002ce245ce, 64'h39724915d70017fd, 64'h1b9ae81222},{64'hc000000, 64'hb080000000000004, 64'he38a5b6d74d6220c, 64'h1f5cd00d960516e5, 64'h3d46b8f51ae993d1, 64'h8f8cc465e},{64'h30000, 64'h5c1a0a0000000000, 64'hb60f9e1776a13165, 64'h9cb99a1e2c428, 64'h70d2a5730, 64'h16b8003720},{64'h0, 64'hb017800000002000, 64'h10bceb61895844, 64'h906d4240d1822044, 64'h1dc388570c000110, 64'he8dc95af4},{64'h4000400000, 64'h615800000000000, 64'h1f516ceb0b3a4c4d, 64'h23d30a1e800464, 64'h1460003a6449c24, 64'h1198001da0},{64'h0, 64'h3017000000004100, 64'h16ba184c3d4305, 64'h3466400021c42000, 64'h1c0869708001990, 64'h32740efe0},{64'hc000000, 64'h7017000000000000, 64'h108c98a101b81d, 64'h89a28000004f8, 64'h74000006a59e8000, 64'h13e8580bc1},{64'h40000, 64'h3014000000003008, 64'hb4aac4c4c9879, 64'haf6797413bf2a144, 64'hf41597d0560a0e81, 64'hebf427395},{64'h2000000000000c0, 64'h4200000000000000, 64'hcfcbb36119b1ee4d, 64'h64a4748e800729, 64'hb7ed1170b59c20, 64'h1a02d670f0},{64'h2000000000, 64'h3000000000000004, 64'h86496be6ea5e480c, 64'h1700a0008e06c6f8, 64'h1d416dc432001196, 64'h15bb8773de},{64'h80000000, 64'h71208e8000000000, 64'he8dd365b50205, 64'h5c3c2a50d8a9000, 64'h3c8480013c0003bc, 64'h1ab2d95ae1},{64'h400003000000000, 64'h7016000000000014, 64'h14d37554b4ca8241, 64'h7923c4314680051a, 64'h143bc006870088ad, 64'h6510c3874},{64'h3000040040, 64'h30f1000000000008, 64'h95ce97b491889, 64'hb7183000bbf12089, 64'h74b796d0622d9d14, 64'h19c1480054},{64'hc01000000000, 64'hf007000000000000, 64'hd4b11510e385b, 64'hc6000001a100018e, 64'h23b001444, 64'h8780021e0},{64'h400000000000002, 64'h3000000000003000, 64'hd53688828c0558a1, 64'h8918430462000515, 64'h10e5b178001403, 64'h8df8a6e40},{64'h300000000000080, 64'h3000000000000000, 64'hb515266e941a105, 64'h17678141a1800663, 64'h49ab704686878906, 64'h1a921f5a6d},{64'h4000000, 64'h4025000000003000, 64'h5a4f8a5135baf493, 64'h6a5001b38006d0, 64'h1cb394734000000, 64'h1ca56a45e0},{64'h2000000000, 64'h7015000000003000, 64'hda31d600af812, 64'h251c00147064000, 64'h59b2b3609acd9aaf, 64'h8af945d0e},{64'h10c0, 64'h8200000000000000, 64'h458d8be55a258b53, 64'h9339a65090786dbd, 64'ha1109c738e724e69, 64'h8b8de3966},{64'h40000c000100, 64'he406000000000008, 64'hcc8f5a9b175d2884, 64'hda3bfb69992a6095, 64'hf44800045f0d5aaa, 64'h18138743fd},{64'h1000000000, 64'h30240d8000005010, 64'h95e2359d1f781, 64'h3244c23815e1e094, 64'h7c00000424000556, 64'h1b4722d58},{64'h10a00000, 64'hf0ba800000001000, 64'he11270836c452304, 64'h1a04f59fc20002ee, 64'h3448cf30a4e3cbb9, 64'h1745192d40},{64'h100c02000000000, 64'hb0f0800000000000, 64'h2496c68bbc1561b, 64'h974d13da88096a2, 64'h1c7dd151b0008fc, 64'hdf04f5ae0},{64'h400000000000, 64'h4600000000000000, 64'h158de93b350252, 64'h5cd6d9c0b1f394, 64'he19c80045bce4000, 64'h3c0750461},{64'h200000000000040, 64'h30a0800000000000, 64'h370cabd095da6315, 64'h12144088000045, 64'h1c3d1407c0003f0, 64'h800000000},{64'h100c0, 64'hb000000000000000, 64'h13bd1a8102181b, 64'h6a4b7546400087, 64'h350437020016e8, 64'h119ec406a0},{64'h30000, 64'hb017000000000000, 64'h104ce4c10db802, 64'hcf665e0422742000, 64'h9dc0b7f6880853d1, 64'h13e85e3a26},{64'h100, 64'h14012380000008, 64'ha04c6ce2b555ee00, 64'h14080038b, 64'h9934000146001060, 64'h14a265178},{64'h860004000000, 64'hb000000000000000, 64'ha9d465d305891803, 64'h3a144d701135c0, 64'he8beed3057d0a000, 64'h5ac3},{64'h300000000010000, 64'h2000, 64'h71535d697b29a000, 64'h8d3a67408edd0592, 64'h35cf5d371a0010cb, 64'h1a05b05bce},{64'hc00000000000, 64'h8408000000000004, 64'h1dce5c669ab6f255, 64'h2dc0010f2d838a, 64'h403c0000f1154b70, 64'h3995570fa},{64'h100, 64'hb02a06a00000000c, 64'h59974320992df81d, 64'h672f232854d1d0b3, 64'h8600023c000849, 64'h5c9606ad0},{64'h20040, 64'h39000000004000, 64'hce574c6a870a7864, 64'h64a0008f5b051b, 64'h8e9ca394000000, 64'h1b9cb71700},{64'h2014000000, 64'h4600000000004000, 64'h4e0dabaf20895862, 64'h4f52a8549712e2, 64'hbcb7cc86840008ec, 64'h196c9f684c},{64'h40000000c0, 64'h6800000001008, 64'h8995bda899a96e00, 64'hc218ae2490204685, 64'hb91280050400054c, 64'h1aaf736ab9},{64'h4000000000, 64'h4018800000000000, 64'h86ccaddcb152439a, 64'h43c0019280067e, 64'hea80000000083c, 64'ha20},{64'h4000020000, 64'hc000000000000004, 64'hc2602ac5a8395, 64'ha96f4079a1c1e712, 64'h70bd8002f8078e9c, 64'h6a5e},{64'h10430000, 64'h3000000000000000, 64'h56937d59172e41b1, 64'h709d57aae8a4fa, 64'h1cb56f0ca19c000, 64'h2de0},{64'h40000000c010000, 64'hf000000000000008, 64'habb6a4c05d8b3, 64'h545d1001474de51a, 64'h513ed9466d001470, 64'h72d6},{64'h40000c000000, 64'h7000000000002000, 64'h168c02b00ab80b, 64'h1f39b59d99344688, 64'h1bf80038fd541a8, 64'h8bc0070e0},{64'h4000080, 64'h3000000000000000, 64'h21558d94c03e63a4, 64'hf45b524000000665, 64'h1cf8002320008c8, 64'h1442675100},{64'h1010001140, 64'h3000000000000000, 64'h84a9d184ee361, 64'h1c00b5dd13632a39, 64'h862e35c6af9745, 64'h298000000},{64'h190000040, 64'h3029800000000000, 64'h8ccd7b868c449861, 64'h8da13e811928d709, 64'h883b9742e853c8d6, 64'h147054014e},{64'h301000008000002, 64'h16a0000000000000, 64'hd4754a1af7519799, 64'h3a3425a190e013, 64'h16bc00005c819c8, 64'h3720},{64'h41800, 64'hb000000000002004, 64'h16d59e284c01f012, 64'h51ba00018f878bc, 64'hfc000006738ad162, 64'he5c5f0f11},{64'h400000000000, 64'hb000000000003008, 64'h16ba5f18097804, 64'h5889e8886dd664, 64'he0000002291e03a8, 64'h224364671},{64'h100000000000000, 64'hf000000000002000, 64'hb83ec9182550c, 64'h5bbb6012800000, 64'h1abc005cce04000, 64'h22f435ac0},{64'h4000000000, 64'h3007800000000004, 64'h13261341389851, 64'h52000000004d0, 64'h351300000000169c, 64'h118a823a38},{64'h418002000000000, 64'h9200000000000004, 64'h44c826052c056c05, 64'h5500147d173503, 64'h1917d7faea52c15c, 64'h300044d0},{64'h800000000040, 64'hb000000000000000, 64'hf957b913582970c, 64'hdd71ade889d105c1, 64'h3dcb0675ad74c8a0, 64'h2284472ca},{64'h300000010010000, 64'hd027c80000000000, 64'hb6e2b182a6c4d, 64'h443770e872d000, 64'had6f5e0000001c6c, 64'he80003a06},{64'h6001400004000080, 64'h7000000000000010, 64'hb8c85aaa4c34b899, 64'hd42ddd5971ac2521, 64'h5e3c57e121588bf8, 64'hb3800605d},{64'h40000c000080, 64'h3000000000000010, 64'hd8c295ba1e099, 64'hb8219475c800023d, 64'ha00000023d6c4e50, 64'h43fc},{64'h1000008000000, 64'h4600000000001000, 64'hba807c284c05789c, 64'heb23fcd0ba1532e8, 64'hcda104e71f72a552, 64'h19d5192343},{64'h0, 64'hc418000000000000, 64'hb176c52b552b664, 64'h40a9c1c48002e3, 64'h1bf82c44a000000, 64'h0},{64'h1000000080, 64'hf000000000000010, 64'hd45460dd2034970c, 64'h2f442cf99fb18241, 64'h40ed8003aa8bd415, 64'h1179da0471},{64'h0, 64'hc207000000003008, 64'h8b098b275a224fba, 64'h2dc554b702103c, 64'hf56b3455ac8a5a28, 64'h10fdf1681d},{64'h200404000000000, 64'hf0e658000000000c, 64'hdac1e9bca7412, 64'hea0960000f400514, 64'h51ce7572f9ba9c0e, 64'h33000715a},{64'h1003000000184, 64'h701b000000000014, 64'ha3af94448c34d859, 64'hc950009d4025c4f5, 64'h60b7f484fb24141d, 64'hd49d70bd7},{64'h2000000000000c0, 64'h200000000000000, 64'hb70d9e255a25eb8a, 64'h8750e98945000397, 64'h2c8dc004fa001476, 64'h16f2bd040a},{64'h2004000000, 64'hb000000000003000, 64'hc9d74a233951cb02, 64'h9470f73400000689, 64'h44cab69122e51ab7, 64'h199f406807},{64'hc01000000100, 64'h27000000000000, 64'h850f6c53754d8b00, 64'he66aca211324c433, 64'h140000073f4308ce, 64'h511a},{64'h20004000100, 64'hf037800000005100, 64'h478bace25c4898a5, 64'hfa51b47cfe80043d, 64'h78c00a55c7ec7471, 64'h16cd1d9961},{64'h400000040080, 64'ha60000000000000c, 64'h43948e18dc4178ba, 64'h36672430bcc00467, 64'h31a88002e9d44838, 64'h1477217454},{64'h10000200c000000, 64'hb800000000000, 64'hc8bd709893200, 64'h739745105800240, 64'h1a24004581719cd, 64'h0},{64'h200000010000000, 64'h4600000000000000, 64'h53d6261d4081f89c, 64'he2191b88000005ba, 64'h119ec52e8ae59a2, 64'h2fd754fa0},{64'h600100200c0, 64'hb018000000000000, 64'hd0d17cdd7489b61a, 64'hbd1853796eed875d, 64'h1a2d60f1d5e8d2, 64'h8bae35c60},{64'h80, 64'ha8da000000000, 64'h8cc98a91385d8100, 64'h7c0fe2cd068005cd, 64'h91987844c1e1349, 64'hbe000462a},{64'h200000004000000, 64'h1cf6814000003000, 64'hb8089c592b8e0b15, 64'ha8057cb1950002e2, 64'h1134061f6b909ca, 64'h14151465a0},{64'h6000000000000080, 64'hd0800000000004, 64'h1113a2af1789c9b4, 64'h9e5b44608c11a227, 64'h968bb4a5bca9c77a, 64'h7134900db},{64'h200000080000000, 64'hdc3b800000000000, 64'hac98b588ace1493, 64'h1485603dc780f65c, 64'h41cb45e0bc03d47d, 64'h1c8053054e},{64'h6200000000000000, 64'hae1b000000000000, 64'h44937d5a97228b92, 64'hd83b0cc59500057c, 64'h7af0f325c63c88a1, 64'h1720873a17},{64'h100030040, 64'h9000000000000000, 64'hb413a362995df075, 64'h67b946adabdd05c7, 64'h559f00067cb44bfd, 64'hd92cf3a0c},{64'h100000008000100, 64'h240000000000000c, 64'h5f174bd8b72a7502, 64'h196755acbe3462ef, 64'h81c8f472de4e0e55, 64'h7a83623d2},{64'hc00000000080, 64'h200000000000010, 64'he2554b68bbcdee8a, 64'h84662ca9d48022e9, 64'hc81e3aa68511575f, 64'h23000015c},{64'h44, 64'h400000000000000c, 64'hb34ab5ec44a6bbc, 64'h912e60851aa9244d, 64'hbda298b294d14b9a, 64'h11b9e75078},{64'h100c0, 64'ha425800000000000, 64'h5b914d68d4326f83, 64'h40ad159ff456af, 64'hedd56456590b38, 64'h130002ce0},{64'h200c0, 64'h8200000000000000, 64'heb934554f809b774, 64'h634000b773f739, 64'hfc263964fa001a2c, 64'h6fac},{64'h10600000, 64'h8400000000001000, 64'h5f4b9540cc3558bb, 64'h79703a56be8002ee, 64'hd2e80066c2c5755, 64'h147c00674c},{64'h6000000000010000, 64'h3000000000000008, 64'h89947ddcb546d80b, 64'hd944c76540420514, 64'h2e4c399691e65091, 64'h1ae8003b17},{64'h4000000, 64'h702b000000000180, 64'hd43e2c9ca171d, 64'h50f73db4800352, 64'hea800720000000, 64'h16f745f220},{64'h10a00000, 64'h5400000000000004, 64'h890c262761029871, 64'h213a7e362f0000b2, 64'h7c00000442001ca6, 64'h112a016811},{64'hc00000011000, 64'h7000000000000000, 64'h8d174a296589d814, 64'h7251130973756c32, 64'h19c31444f4790f0, 64'h10fa356700},{64'h8000000, 64'hc600000000001000, 64'ha2178a616429ac7c, 64'h7051fb9973084072, 64'h10ff445218211442, 64'hc0c3708a2},{64'h8000000, 64'h714985c000000000, 64'h11508ddebaaacd02, 64'h673a1c22842238, 64'h1440006a3000000, 64'hc08004c60},{64'h218001010000000, 64'h3000000000000000, 64'h7614ade6a602d841, 64'h21155ce59c889572, 64'h282fd15a43001167, 64'hecba17440},{64'h3000000080, 64'hb000000000001000, 64'h6a495aaf544e3405, 64'h5c57248a0005bb, 64'h2c8d000228409abc, 64'hbaebe2007},{64'h804000000000, 64'h7000000000000000, 64'h5d0e7d2775b14102, 64'h510978bc8006ae, 64'haa0006895f0eac, 64'hbaa875c70},{64'h1060000000142, 64'h3000000000000008, 64'h8ce99caec43e80b1, 64'h4ea0314632c03d, 64'hd53980c5ad89a060, 64'h5059},{64'h460000000000, 64'ha800000004100, 64'h14506cd6c9509800, 64'h5250492d6e0004fc, 64'h495e1d85c95d6ea8, 64'h145d14bb01},{64'h11000, 64'h600000000000000, 64'h3ecbbc5506da72a3, 64'h5751e14c8d51881e, 64'h1a5790762a41480, 64'h81142280},{64'h4000000000c0, 64'hd1580800000008, 64'hb8cf8c13753a7200, 64'h73400007d18057, 64'ha9618f30bd001cd0, 64'h898f0721d},{64'h4004000000, 64'h4400000000000000, 64'h5cd05caa9c5d8343, 64'h263b1c55aa02b056, 64'h19960e44c5d448e, 64'h16880029c0},{64'h40000c041000, 64'h316a810000000000, 64'h1753dcd88678a1, 64'hd63955b4865d0daa, 64'h194134667d530192, 64'h1352cf504d},{64'h40, 64'hc40000000000000c, 64'hdf164c5706a90c9b, 64'h8a00d988402f9, 64'h29a3f9c738000000, 64'h196baa235e},{64'h400000000000000, 64'hc0b1800000003000, 64'hb74dbba8814aa14c, 64'h394000e52c5294, 64'h87c22000000d90, 64'h1c56de0000},{64'h80000c000000, 64'h7000000000001000, 64'h352852f548ed813, 64'h2e784149420708, 64'hb3b4268be1d160, 64'h11bc2c0580},{64'h40080, 64'h3016000000000000, 64'h1309aaad77c26369, 64'h23814d9a745add, 64'h8785f54c178000, 64'h1d811d0000},{64'hc00014200080, 64'hb000000000000010, 64'h9f8f9b64c486f843, 64'h165adbab9fe4b72d, 64'h24e49a56b10599c0, 64'h18c0165b37},{64'h501000000030004, 64'h7000000000000000, 64'h5e6f4c56d64101bd, 64'h428019416262fb, 64'h7d18f930f1084030, 64'h726d},{64'h400000004000000, 64'h260000000000000c, 64'h5e4a5b6b210df881, 64'h8e3b35e4e8381368, 64'h90036a4733755c83, 64'h14e00068ba},{64'h2000000000, 64'h717981e000004000, 64'hb436960c22315, 64'h100000000000662, 64'h668001cb6, 64'h22c006840},{64'h400000000000080, 64'h3000000000000184, 64'hb98e26011c2898b1, 64'he63b021d8a21e6ad, 64'h6597c063b2e7c8fa, 64'h112f578bfb},{64'h200000000000000, 64'h303806a000000000, 64'hc8cf6e2537457715, 64'h8438a000ab33f2dc, 64'h599c7560000001d0, 64'h11ad6f680d},{64'h200003000000000, 64'h3018800000000000, 64'ha18b936b755a8914, 64'h674ba00171286511, 64'hd422c005c8ae9ac6, 64'h11a8735108},{64'hc02000000000, 64'h4200000000000000, 64'h5f084aeb2bd1ee54, 64'h2fa7645009808b, 64'h452ea305bac90c, 64'h228000000},{64'h3000020000, 64'h1000, 64'h1662f49350f00, 64'h2280019cdb6394, 64'h687f107000001724, 64'hece317454},{64'h10000000000c0, 64'h4000000000000000, 64'hb6092616c15aa193, 64'h376a2000000005c9, 64'h45f985a88, 64'h16c80050e0},{64'h2000000000, 64'h3000000000001180, 64'h3108c94f00ef81a, 64'h7f01694805a7a518, 64'h13aa730169fcbe6, 64'hbaf58cf40},{64'h0, 64'h2b059700000000, 64'he2cf9c54dac9d400, 64'h19e281c0005b8, 64'h3029000072001300, 64'h14083957ae},{64'h100000000000000, 64'h406000000000000, 64'h2c49a3af35d94344, 64'h1460002fa, 64'hec57f000000330, 64'h1478580000},{64'h2000000000000000, 64'h7000000000000010, 64'hb16bb5101509802, 64'h2c6d409c00000466, 64'h531896c2d8001484, 64'h11a1405174},{64'h3000200000, 64'hb000000000002000, 64'he64d4ba33bd98804, 64'h73546bcca8f6a8, 64'h3c87b610ce0008a4, 64'h1725752b2a},{64'h200001000000000, 64'h600000000000000, 64'hb7568dba540b3, 64'h4681c0b6a34000, 64'h59a054d5a6001134, 64'h66b},{64'h110000000000000, 64'h8000000000000000, 64'h929d68d185585b, 64'h5d00400000000662, 64'h1a3682f32001743, 64'h1978030000},{64'h300000014040000, 64'h4000000000002000, 64'h1a97926c80c09874, 64'h3a2190997374566c, 64'h29d54fe4740008a2, 64'h23737228c},{64'h2000000000, 64'hc600000000001000, 64'hebc6cb4a9b0ac, 64'h12458430e57546f8, 64'hd1cb171684e58bae, 64'h16f7552e22},{64'h400000000000, 64'h4437000000000000, 64'he1ca5b5967d66994, 64'hd60008e3a3000, 64'h7c3580170f02c000, 64'h35b880591},{64'hc00000020000, 64'hda1a016000000000, 64'h7959e2ef4b112b4, 64'h87670059755a5630, 64'h1c28005bfe1dc33, 64'h6d60},{64'h100c00000000000, 64'h7130000000000000, 64'hcbc60a7cac20d, 64'h264204840335f180, 64'he4d20507e4c0b6, 64'h1488665220},{64'h400000000c000000, 64'h5f41800000000010, 64'he5c84a9b69c64105, 64'hda70db11a3a0, 64'h1fc9c0e234408000, 64'h1cc00065bd},{64'hc00000000000, 64'hf000000000000008, 64'he7d6ed45a8104, 64'hf038df408000000, 64'h15277d72f06d9a0, 64'h1990007230},{64'h400000008000140, 64'h70080d0000006080, 64'h88cf2c9e6c4e986c, 64'hf7685b991180001f, 64'h95c86db55c444889, 64'h8627db63},{64'h300400000000000, 64'h29800000000000, 64'hf5c291ba9cd00, 64'h678e44e2b9108a, 64'h359d4433b3c11cfc, 64'h6ac0},{64'h1400000000100, 64'hf000000000002004, 64'hb8935d6cd1aa9893, 64'h520cf54819e057, 64'hf5ab70c5a31659e8, 64'hb7da2681a},{64'h300000000000040, 64'hc400000000000000, 64'hb849ae20d9c9f4ba, 64'hb0000001752e150d, 64'hf54440009a76448a, 64'h19eb0846bc},{64'h4000000, 64'h10, 64'h158dd095d1c27c, 64'h502fba14e5000368, 64'hc48122a2348a942a, 64'hfc8007158},{64'h30000, 64'h8405800000000000, 64'h5c8d43e119b981a5, 64'h8a57250c, 64'hb1440004d8084a08, 64'h168004bc0},{64'h300004000000000, 64'h8200000000000008, 64'hced585d6f4595863, 64'h366a39dd1b000016, 64'hd5ac4004f41e0b3c, 64'h633c6b18},{64'h20000, 64'h81584000000000, 64'h178a56fa3a6100, 64'h71600005c00000, 64'h20b913d4c25c93fc, 64'h16f38c502b},{64'h0, 64'h8200000000000000, 64'ha08c6bd4e1a1624c, 64'h702fa2a8cda54518, 64'h1800000073001412, 64'he4286390a},{64'h3004000000, 64'hc02b000000000000, 64'h108dd14526ab94, 64'h6c51f501c0800000, 64'he4000002f80e5495, 64'h3b00},{64'h3014000102, 64'h30f5800000002000, 64'hb2e26145c02711d, 64'h673abd551c0002f3, 64'he9478682d9d55ce5, 64'h11a55b2ea1},{64'h46, 64'h4000000000000000, 64'hd5745e1f19a92263, 64'hce4fe73819800733, 64'h12999d5a20013f9, 64'h16b0000000},{64'h440010000000, 64'h8600000000005000, 64'h709064a2d98a9843, 64'h23fba11a761732, 64'h19c02dfd1a000, 64'h10ff320000},{64'h40000, 64'h148a6c00000000, 64'h176e2d51800000, 64'h58474d444270a000, 64'hdc8a00000000035b, 64'h1c38200c},{64'h0, 64'h2400000000001180, 64'h134c58a106ab04, 64'h234282d1160002da, 64'h9c000002de7d11d6, 64'h19bf46a9c8},{64'h400000000000, 64'hf000000000002000, 64'he8d17aeca7524304, 64'h5c8d340134d556, 64'h4b8fa472d1ac0f8, 64'h1aac015c20},{64'h0, 64'h3489e000001000, 64'hdb575e270aaad26d, 64'h70c0219c851646, 64'h14b000010000000, 64'h1c440952c0},{64'h300000000000000, 64'hc200000000000000, 64'haab26e4d2c295, 64'h9300000000000056, 64'h1ce5f886c0001c3f, 64'h90b46196d},{64'hc00014000184, 64'hb000000000004000, 64'h89a9b2c6e8a14169, 64'h74eb46829068019, 64'h4c8391b727a11421, 64'h146c005231},{64'h4000030000, 64'h1600000000001008, 64'h138b5f584d80a1, 64'h1b6ac5d5524106ac, 64'hba95d3b4624294, 64'h1cc61f3a30},{64'h20040, 64'h4000000000003000, 64'he7e18d9c9368d, 64'h662228a5bece5039, 64'hb4000005b67d1490, 64'h1bf6af5228},{64'h200000000000040, 64'h6400000000000000, 64'h6e137ad518092e05, 64'hd3330001951c7447, 64'h456df5639600088d, 64'h231d16807},{64'h0, 64'h614000000000000, 64'h7355939375b62255, 64'h1cc661c8c0022e, 64'hd11a13a2000000, 64'h1721185900},{64'h4020000, 64'h4000000000000000, 64'h179bad24a14363, 64'h67b765484980da, 64'hec8b23b22c334000, 64'he719939c8},{64'h800000000000, 64'h4600000000000004, 64'h6e0bb358f7212a9d, 64'h67ab79860bb5c3, 64'hd6f2cc5d7d00000, 64'he58c367b3},{64'h2004000000, 64'hc600000000000000, 64'h8a49aad8d9ca8f45, 64'h50be71149f4058, 64'h137344455a208d4, 64'h1cc00f0000},{64'h4000020000, 64'h301b000000000000, 64'ha2084ce95bbd8369, 64'h4eaa15446342e5, 64'h13d000000001a14, 64'h1ba510e20},{64'h500000000000000, 64'h3000000000004000, 64'h16534dd921554102, 64'h3672a00148374520, 64'h2fe824d88d9caa, 64'h8ef3cbd20},{64'h40010000000, 64'h820000000000000c, 64'h88cf54615952f66b, 64'h2d000bc8002f2, 64'he0000002e5b7bcf8, 64'h1120007197},{64'h4300000000040000, 64'h3000000000000004, 64'hbc575a074c0ed881, 64'h37070cd403735505, 64'h1abfdd8242000be0, 64'h8eaf2391a},{64'hc02000000000, 64'h805a000000000, 64'h138d6f24b91800, 64'h51e000000000f8, 64'hf4ba80073b000b64, 64'h1468002ba1},{64'h1400004000100, 64'hb000000000000000, 64'h8e2c50a481817805, 64'h6ab718e3000669, 64'h316b38c665b79740, 64'h16509c5bce},{64'h2000200100, 64'hd58d8000000000, 64'ha0934d1487c09800, 64'h4ff73b413315cd, 64'hb4e43323389d5a34, 64'he1800390c},{64'h400000000000, 64'h4000000000000, 64'h94d55b68fba9cc00, 64'h6849fd1d27f668, 64'h81342739450000, 64'hd80},{64'hc000000, 64'ha800000000000008, 64'h2093bd5b693d811a, 64'h22475141132145b2, 64'h6400000444001ac6, 64'hb7ada66f5},{64'h30080, 64'h4000000000000000, 64'h8cd69a5d78a161a5, 64'hbac01459, 64'h19b800616ce8000, 64'h19d32866e0},{64'h1003008010000, 64'h7000000000000000, 64'h14484bd4e65c9805, 64'hec5c92dda6f25672, 64'h58200b7463bb1d26, 64'h1d24b752ea},{64'hc00000000000, 64'hd400000000001000, 64'hd4cdec8daa25d, 64'h2123e0ed758005d6, 64'h14b43470f001a31, 64'h4f880000},{64'h1000000140, 64'h600000000004000, 64'h41149da0d0464249, 64'h1a70ee0404000017, 64'h34b87000001c9d, 64'h640920a0},{64'h1000000000, 64'h809a00000000000c, 64'hd80d9ca37105988a, 64'h9351e0009e81c038, 64'h9c938b62e4e59427, 64'ha74},{64'hc000004, 64'h361d46000000010, 64'hd5ab6b2377c89875, 64'hf9039abc420693b5, 64'hf93f0004542156d9, 64'h4280051b9},{64'h104100c000000, 64'h4000000000000000, 64'hbab11478a7074, 64'h6c2235bdcf80073e, 64'h5a0008073b6f495, 64'he59b965a5},{64'h800000000000, 64'h8600000000000004, 64'he6d46da2b9a12062, 64'h39cb90ceb9b5c2, 64'h90000006ad689b98, 64'h1652b13a3b},{64'h0, 64'h37800000001000, 64'h149585ec99ad0295, 64'hd53aa0000000019a, 64'h1ac1, 64'h8c4000a60},{64'h4600400000050000, 64'hb0ab800000003010, 64'h5f81b6204c0e381c, 64'h4504c574628102, 64'h3a01e3ba2d2f0000, 64'hedd7f6657},{64'h6000800004000000, 64'h0, 64'hdb179a656a81f800, 64'h5bd4448a394398, 64'h2e730006819c1440, 64'he689b1877},{64'h3000000040, 64'hc400000000000000, 64'h1ad5be2c944d9483, 64'h7a73900000000453, 64'h12a86c462cc9a26, 64'h50c0},{64'h400003014020000, 64'hf018800000000000, 64'h5a8a602e5689d81b, 64'hd70011b795304, 64'hd400e6e504dd5a04, 64'hc196b13a2},{64'h4000080, 64'hea00000000000000, 64'hde175a6ca439a30b, 64'h4472be71c337a521, 64'hb1051d270ed111b7, 64'h1160947388},{64'h403008000000, 64'hdd17800000000000, 64'hbc4d4e10c5aab3a5, 64'h82ff0001c0005e4, 64'hf41c8002ffd01d07, 64'h1124385e4c},{64'h1000, 64'h2c00000000001000, 64'hb8bc09c058abd, 64'h720019ad21d20, 64'h11785f45e0e5490, 64'h17943a0000},{64'h3000011000, 64'hb000000000000000, 64'hd5527a6cd8099813, 64'h9c5d000147e39a38, 64'h556f0002eb0011cc, 64'h1aa91d598d},{64'h0, 64'h7029000000000000, 64'h484dd165b14104, 64'h173ce74e36e8662, 64'h8005d6001758, 64'h700065e0},{64'h200000000000040, 64'h8000000000000010, 64'he41344a2cbbab0b2, 64'h2268e0003638f505, 64'hb0e46ec6840f9a38, 64'h1c880008db},{64'h2000001800, 64'h3017000000000000, 64'h108c96f6dea81d, 64'h3f00013fe3a800, 64'h44000001060008a4, 64'hada242de1},{64'h1000000000, 64'hf000000000000000, 64'ha08a40932185d802, 64'h3646c7a53f800616, 64'h4951116, 64'h16d6340000},{64'h100000000000000, 64'hb02480000000000c, 64'he6919ca8fb86c01b, 64'h2036d64e, 64'h19be9616e000290, 64'h19d39c7490},{64'h1000000000, 64'h607000000004000, 64'h1317aa516106986c, 64'h2544a74c90aec5d8, 64'h5d4b35652c149766, 64'h16f8a410d},{64'h8000000, 64'hed410d2000000004, 64'h9e8d9ae2a931eead, 64'h243768ed2365d7, 64'h9d1880031a000000, 64'h8c00068f3},{64'h300000000000000, 64'hf000000000002000, 64'h2d956626ea216115, 64'h4870fd21478332e4, 64'h8dc0024ee85d0b, 64'h144d4271a0},{64'h400000000000, 64'hdc2a000000000000, 64'hd1acdea8592305, 64'h92742e4801ba1452, 64'h93df572d07801b, 64'h1c700010a0},{64'h1402010000000, 64'h4615000000000000, 64'h2117ce48ad217b3, 64'hdf2f9d55aa977338, 64'h13f5c83b177d6dd, 64'h438000000},{64'h4000006, 64'hf000000000000000, 64'hd02f44675a36c205, 64'h992dfe300000073f, 64'h39722cc000001c61, 64'h5987},{64'h400005000000000, 64'h4200000000000000, 64'hc50a049ae2363, 64'h586680019a000737, 64'h1c64003b0cc96b7, 64'h0},{64'h1000004000000, 64'hf000000000000008, 64'hd34270c32c06988b, 64'h6b15bda6800235, 64'h80b795d3872088d0, 64'h8d9053b70},{64'h10080, 64'hf000000000000000, 64'h41104a28bbb1b30b, 64'h9b2fe5f114400187, 64'h13f06a2fe0008a0, 64'hbfc000000},{64'hc000000, 64'h7000000000000080, 64'h98ce9c98dc42e20c, 64'hb7511b79440c2184, 64'h1408004eaa056d8, 64'h1cb5cdd600},{64'h6100000000000000, 64'h8000000000000008, 64'he50cbbeb1b4153a3, 64'h16a001b680072a, 64'h6364004e0001410, 64'h1bb39646fd},{64'h30000, 64'h2c00000000000080, 64'h5dd7a260e102581a, 64'hae6aa3cdcaf7a70c, 64'he81193a0001ab1, 64'hb5d83a320},{64'h400000, 64'h4600000000000004, 64'hd5cc8b9536caf0b5, 64'h3a5e7200000072, 64'h61790006640016b0, 64'h1a0328459d},{64'h10000000c0, 64'hb000000000004008, 64'h35782d0900acc0b, 64'h9872ee581cb915e5, 64'h34000000180019d7, 64'h4e8d5e5a},{64'h300001000050100, 64'ha20a000000002000, 64'h7795bcc29c057893, 64'h1123e2100e5de039, 64'h11d46c386045494, 64'h11d46c0220},{64'h803000000000, 64'hb0d4800000000004, 64'hd1cf546b3b86581b, 64'hf2002e101d0006ab, 64'h78128005bdbc8e5e, 64'h1993486abe},{64'h2000000000, 64'h190d0000000000, 64'hfa46ec4ae6000, 64'h47044e700000007c, 64'hc9ce00000000175f, 64'hbfb7d2fe4},{64'h100004000000000, 64'hb000000000002180, 64'hc4cd0b506d88c, 64'h68fe61cc338670, 64'h7d7656f03ac6cd14, 64'h1c8e3daba8},{64'h2200000000030000, 64'hf000000000000010, 64'h72557da6ea354012, 64'h456ce96f5c9658, 64'h9f13f3a358001158, 64'h10332d0a78},{64'h40, 64'h840000000000000c, 64'hbacd4ce08955d76d, 64'h2246da584e800505, 64'hc1e00069c001a70, 64'h2a18374d6},{64'h0, 64'h600000000000004, 64'he8c1345dd829a, 64'h112a0844c, 64'h9d0b89f38660cc18, 64'h1ce7566758},{64'h8000040400c0, 64'h6800000000000000, 64'he6cf6c2cc5a5c00d, 64'h44b4253d4f55d9, 64'h4c8985352d000298, 64'h1ce3742261},{64'hc011000, 64'hf000000000000000, 64'h49cd5c15565d2814, 64'hb7513e34ed51ac6d, 64'h1a00016c000938, 64'h24e0},{64'hc04080400000, 64'hae00000000000000, 64'hc019e00cc0e3053, 64'ha1e915d71621403c, 64'hbdc8b9024f001a27, 64'h23910080},{64'h10080, 64'hb0a1204000000000, 64'he8175e12d652a305, 64'h972521dd0c06007, 64'h8800000000000dd8, 64'h396e},{64'h10000, 64'hf000000000003000, 64'h17aad5010e3804, 64'h4468e001aaece000, 64'h8da38005d6d20eff, 64'h1d040068e0},{64'h40004000100, 64'h3000000000000000, 64'hcd125bd51602a371, 64'h75719d613d2825d1, 64'h6dabb6e5c9747aba, 64'h1cd800506e},{64'h10080, 64'hc600000000000000, 64'h86aeb1532909d, 64'h234001ac4206b1, 64'h1a20003b741cb78, 64'h1a70002c40},{64'h300000010000040, 64'h5000000000000000, 64'h9e8c2620a149e00d, 64'h685e31c600069b, 64'h116c6d386744368, 64'he89b90da0},{64'h3000020000, 64'hf149800000001000, 64'h910d5410978dd80d, 64'h2ffa208a6ce5c8, 64'h1722925bcb30e8c, 64'h141e735240},{64'h40, 64'h4400000000000010, 64'habb58fb4d2375, 64'h2ce0005b8c2185, 64'h503001bb0, 64'h5c0004690},{64'h102200c0, 64'h3000000000000000, 64'hcf838028440a58a9, 64'h6416fa0ab7f3e72b, 64'h1cf31950200140a, 64'h1c3b7d0000},{64'h508002000040000, 64'h7000000000000000, 64'h8e8e8c2adba12361, 64'h2a5ac5d490d5f6ae, 64'h1c5519ba15d5ab7, 64'h11d86d6800},{64'h6200000000000000, 64'hb000000000000000, 64'h174a1f59aa21b4, 64'h120000000072e, 64'hef7940901c000000, 64'h48006b1c},{64'h200100, 64'h0, 64'h5d4d44824159c300, 64'h9672da4a4281151f, 64'h429752baa5842a, 64'hef8530000},{64'h201000000000040, 64'h295000000000000c, 64'ha08f4c5aeb858881, 64'h565045f1aa8003bd, 64'h29aaf9e10b0ec08f, 64'h139800399e},{64'h0, 64'hf000000000001000, 64'hd5549c648bb56203, 64'h72ce50908005d8, 64'hb1aa80009ae71794, 64'h1a44006fed},{64'h30000, 64'h8000000000000004, 64'h3dd35c994bd9c27a, 64'h46c465a3d1903a, 64'hdcf6000000000000, 64'h19cb1c2ff8},{64'h800000010006, 64'h5000000000000000, 64'h89f3bd64c586d802, 64'h6545fdcc534671, 64'hfc000002df001950, 64'he51ad6745},{64'h4000080, 64'h8000000000000000, 64'hbacd501892854, 64'h457b8d60800393, 64'h4cc180013ca59718, 64'h461},{64'h8000000, 64'hc600000000000004, 64'ha1d0a4c2e601587a, 64'h5d98654380013e, 64'h6ac761a74, 64'h113a663070},{64'h30000, 64'hb000000000000000, 64'h144dd130b9e205, 64'h57e54112d0c234, 64'hb8000002263d8c1c, 64'h16e96e5ba5},{64'h100000000000000, 64'h4600000000002000, 64'h892933585eeb5, 64'h8e042001d0825000, 64'h3889f4e00000029f, 64'h1ce748170d},{64'h20000000c0, 64'hb000000000000000, 64'h8b0b93691026a112, 64'h742e860ca918324f, 64'h810b81202400093d, 64'h90007222},{64'h30000, 64'h415000000000000, 64'h73cd43a6bac692bb, 64'h11063045cb5cf37a, 64'h14e59aa07414c298, 64'h741},{64'h4000c00000000000, 64'h3138c1e000004000, 64'h63556dd960a88e59, 64'hed0d8bb4ed0003b4, 64'h82000003c11b175a, 64'h1d69c745e},{64'h408000008000000, 64'h38000000000000, 64'h30914ce97b3c9200, 64'h5c9a0800000186, 64'he036747e91e89c88, 64'h60004e62},{64'h500c02000000100, 64'h3000000000000000, 64'ha590462ebb4d4179, 64'h5e40ec2a2f2003, 64'hd1995196b3d11abc, 64'h14b8007373},{64'h4000000, 64'h7800000003000, 64'hd597a2253ab56200, 64'he42dfb911280044a, 64'h45178000da824dda, 64'h1a77573a2b},{64'hc000000, 64'h207000000000008, 64'h576268fb457354, 64'h5075bcaf80059c, 64'ha4010c45c85bc000, 64'h11293a54},{64'hc000080, 64'h8200000000000000, 64'h2dc96ad1763e9375, 64'ha05bd744b50ac511, 64'h294956a3a0450813, 64'hd79157400},{64'h300800000000000, 64'h261b800000000000, 64'he10dad14b8be0972, 64'h52c8ad4b3870a6, 64'hfc61c002e18b5030, 64'h1cb40e70ed},{64'h30040, 64'hc400000000000000, 64'hcb174d6707cad452, 64'h750da001cf40067d, 64'h65a000000000140d, 64'h1ac0002c4b},{64'h0, 64'hc600000000000000, 64'hd38cb8a2a0825842, 64'h502d018cb4e67c, 64'h9400000012041408, 64'h11dc247309},{64'h40, 64'hc407000000000000, 64'h57d54de0b95a9353, 64'h10a14dac000525, 64'h1990002eadc1ac0, 64'h1ca80072a0},{64'h0, 64'hf039000000005110, 64'h106510f53ae104, 64'h3a442001abb56156, 64'h57918173ce3d4b4, 64'h25df8096},{64'h180000040, 64'h7000000000000000, 64'hde0bb36b2a39e264, 64'hf3dd805800000505, 64'h5d49000524915ab6, 64'h1ce01708c0},{64'h40, 64'hc600000000000000, 64'h8d899ad8f7494245, 64'h72dc708d0006ab, 64'he51b91b46e1c4848, 64'h468c},{64'h1000, 64'hd600000000003000, 64'h148358f75d411c, 64'h8835a9c08cf9cc4c, 64'h240000044e85cbfa, 64'h19cf2f394a},{64'h400000000000, 64'h4608000000002000, 64'h15167ba3358a4a0a, 64'h3966ec0000052c, 64'hbd77840675084000, 64'he574e396b},{64'h100800000040000, 64'hc600000000000000, 64'h1f4b6b153925f8b5, 64'h5c7e59c67942de, 64'hc1d6f69f574000, 64'h1b6a394720},{64'h400000300c000000, 64'h4, 64'h289ba9afb551300, 64'h137610280000050f, 64'h5eb7151000000c25, 64'h7b80b44fd},{64'h2000803000000000, 64'h0, 64'h11d79a42d6091100, 64'h4a69428cbf8002fe, 64'hbb78000227d208df, 64'h168265bb5},{64'h46, 64'h400000000000000, 64'h4a6cbe229952767a, 64'h810246045038c743, 64'hc1a77a1000000091, 64'h1d7e1c7442},{64'h8010000, 64'h710048000000000c, 64'hbb915cdb5506981a, 64'h722e9e6cc1eee5bc, 64'hfc1d2de025b31cdb, 64'h45b0},{64'h403000000000, 64'h26000000000000, 64'hbb555de119b5f600, 64'h6c538a800000039f, 64'he16eac03971d022c, 64'h1772385ba8},{64'h40040, 64'hb028800000000000, 64'ha0897aef3429ac04, 64'h5dbe8808cc33b5, 64'h13e9236ae48d3b8, 64'h200018a0},{64'h0, 64'h61a800000000000, 64'hd53dccc5e029a, 64'h8cb6e738, 64'h1e0001f0155cbc, 64'h7360},{64'h10000, 64'hf000000000000000, 64'h8aada8e1059803, 64'h90000001794023b4, 64'hda58003b60a1699, 64'h14bc006960},{64'hc00008000040, 64'h3000000000000000, 64'he797aad4f65a2e14, 64'h5c9b8c6200044b, 64'h19610033a3e80498, 64'h1abdc60047},{64'h8000000, 64'h3015000000000000, 64'h982eed7cd8305, 64'h6a2df000d500039e, 64'h591dd3ba0008a1, 64'h828972530},{64'h1000000000, 64'h0, 64'hd4bad41c1028b, 64'h8110c00105021042, 64'h89c388610c001d07, 64'h4580},{64'h1000, 64'h200000000000000, 64'h216aadcd9322355, 64'hf05e012dc3e96dcc, 64'h14b856758a5dd62, 64'h6b00},{64'h4000000, 64'h8600000000002000, 64'h119c98d7baf055, 64'h6e2eb0014a064528, 64'h1a623b681d30190, 64'h11e7406500},{64'h3004000000, 64'h8400000000000000, 64'he84d8e1907d2b64a, 64'h805035d00000069d, 64'ha9b95300001cc5, 64'h1b88a60000},{64'h400000000001800, 64'h1a00000000000004, 64'he4c6e4c4d820a, 64'hf3000001ac698eac, 64'h1c8f9045e2b1cf2, 64'h2280072b0},{64'h5010000000, 64'hf000000000000000, 64'h77d068ace0c50303, 64'h8802317d741df5d0, 64'hc0c1700000029c, 64'h14c0005300},{64'h200400010600000, 64'hb0d0000000000000, 64'he9889aab1b8a9815, 64'h415d7e721dba6076, 64'hf177406525bbd778, 64'h11b87202f0},{64'h400000000000, 64'h702400000000000c, 64'ha4956ded45be300a, 64'h7246e0011b80050e, 64'h1c8dc0046fa49330, 64'h124000673d},{64'h10600000, 64'h200000000000008, 64'h128d1e8bac98b4, 64'h53689cea20000000, 64'he580044fd3d4b0, 64'hdf02d3950},{64'h4000000000, 64'h4600000000000000, 64'hdb4c40414c3d2284, 64'h7e6748ed1d800728, 64'h7577e3900000036c, 64'h38000672c},{64'h40, 64'h5a00000000000000, 64'h54534514b95ae204, 64'h8173849c8f9272df, 64'h2c000002dc2e1ce3, 64'h4730},{64'h100002000000000, 64'h30b0000000004000, 64'h137d611906eea1, 64'h4468800000000094, 64'hb74a400000089f, 64'h5c40b8000},{64'h4000080, 64'hb000000000003080, 64'he5826e071c02d81c, 64'h695e88c08b02ff, 64'h1116b7f5e1e59d18, 64'h1a57b1c3e0},{64'h400000, 64'h8600000000000004, 64'he8935c1edb82b462, 64'h3036120483f59c, 64'h5bc000000, 64'h50007450},{64'h10200000, 64'h3000000000000000, 64'hb00eb0a84402b8b9, 64'h13e6ee98005dd, 64'h11c0005ba000000, 64'h3a8005420},{64'h200000000040000, 64'h3000000000001000, 64'h57c2bb82a1810ca1, 64'h8d50299442c002de, 64'h16eddc2de771ab8, 64'h17768b4710},{64'h30000, 64'h4200000000000000, 64'hd8bdd7b4a6282, 64'h736091d151a69c, 64'hc20a2247424000, 64'h1b9b4f3080},{64'h80000c0, 64'h0, 64'h169a54d655e192, 64'h75e7b597229652f, 64'hed8076960002a0, 64'h1480300e0},{64'h100000000000000, 64'hc626012000000000, 64'h824d546b0c050ea4, 64'hb973e01c5c80044a, 64'h1a5ed144e2e5720, 64'h0},{64'h300000010000000, 64'hc200000000000000, 64'h117d2d7741a294, 64'hf72ff6ec00000722, 64'h4494c2201e000898, 64'h1c93af38d7},{64'h30000, 64'h4400000000000000, 64'hd5496e2ce42e6184, 64'h562fe098b5400458, 64'h1cc0103bb85c433, 64'h113b17300},{64'h800000000000, 64'hc618010000000000, 64'h99e14d65e51b3, 64'h9758315780000ac, 64'h2600070f48d4b8, 64'h0},{64'h402000000000, 64'h6400000000003000, 64'hf9e0368019414, 64'h4c5e1ca94c00052e, 64'hcc2f80052f195d67, 64'h1ace956800},{64'h400000000080, 64'he200000000000000, 64'h1665153189e90a, 64'h196e20000d800529, 64'hb1011699e54ba8, 64'hc8004790},{64'h300004014000000, 64'h7000000000001000, 64'h10608727a1b1a1, 64'h80825bcdcf2f7000, 64'h19caf4915ed24095, 64'h1d17574681},{64'h1060000000000, 64'hb140000000000000, 64'hdabd2a0cd621b, 64'h73dbac00000000, 64'h8000000075607178, 64'hf00001121},{64'h800010000040, 64'h3000000000000000, 64'h4841520531817881, 64'hd9bbc030003bf, 64'h83b8b95dd000000, 64'h1e1225311},{64'hc02000000100, 64'h3014000000000000, 64'he9b76a44b98d9805, 64'h84510e1d49000187, 64'h1a3983471e1d77f, 64'h3989f4e60},{64'h0, 64'h3026068000000000, 64'h16cd4e1f19c94302, 64'h3002991be96526, 64'hb8000000a8000c00, 64'h14a0003946},{64'h200000000000000, 64'h8600000000001000, 64'h8ed6ba21392960ab, 64'he0000000006f0, 64'hfda84004720019d0, 64'h1787966641},{64'h418000000000000, 64'hae00000000000000, 64'h9b0a0a08d6e04, 64'h70825d1df87694, 64'h1639f0e774ee8, 64'h5cb4b04e0},{64'h800004000000, 64'h3000000000003000, 64'h76cf9c2ca4ba5502, 64'h73922c93ee65cc, 64'h2ddd61ab8, 64'h905dc5160},{64'h200c00000000000, 64'hb000000000000004, 64'h605053ef348ab815, 64'h70208811000301, 64'h1978c006952c5cb0, 64'h11af06951},{64'h200c0, 64'hee00000000000000, 64'h2495e2934424113, 64'h935bc01cc0fa445b, 64'h169877526165d1e, 64'h11ea3c0000},{64'h80, 64'h1b80000000000c, 64'hd2d59e12d439f193, 64'hdf752b7c008005df, 64'h17982e5e60f9d4a, 64'h1a60497470},{64'h2000000000000c0, 64'h5000000000000004, 64'h77114ce14931eebb, 64'h4f4f4d3c490003a7, 64'h391c4005bb0b4ee3, 64'h1419dd5dd2},{64'hc000040, 64'he000000000000000, 64'h46917cef44a24202, 64'h176af05c000002df, 64'h1bf8253b9e70860, 64'h69e0},{64'h408000000000000, 64'h2600000000000000, 64'h6117809ec181aa89, 64'h460522dd799845e6, 64'hbd8480e475a58, 64'h1a7cab23c0},{64'h860000010000, 64'ha007000000000010, 64'h344f9aa91b553714, 64'h95c82e54be19744, 64'h69698da697b97d00, 64'h113ba346f3},{64'hc00000000000, 64'h4301826000000000, 64'h244bbb6d14c98245, 64'h493c00000000001e, 64'h24800741744f00, 64'he00000920},{64'h0, 64'hb000000000001180, 64'h5bcc5461793d020d, 64'h10d810056, 64'h1a7c002dc548000, 64'h1c9515c5a0},{64'h100002000000000, 64'h7000000000000000, 64'h130e7dd54182d80d, 64'h57697a5c8a0005e0, 64'h1cc400212001ab4, 64'h8a8000140},{64'h8c020000, 64'hb000000000000010, 64'h1472057b06331a, 64'h97f59d3178433144, 64'h55a018430800091e, 64'h196866017a},{64'h3000000000, 64'h5600000000002000, 64'h600db398808eb312, 64'ha92ea0094c7a9752, 64'hb2019304001a64, 64'h14ac000240},{64'h403000000000, 64'h8400000000000000, 64'hbdd78bab3b49806a, 64'hbb8002ee, 64'h1a480072bbe00e4, 64'h0},{64'h300002000010000, 64'hf000000000000000, 64'h2e007e074c0ed865, 64'hb8170001abea30a8, 64'hc14556930017a4, 64'h320555dc0},{64'h20000000c000000, 64'h3000000000000000, 64'h389b3651baaa112, 64'h45f03977842172, 64'h14c63801c0003a8, 64'hf04000000},{64'h4030000, 64'hb000000000000000, 64'hd01375c35a360205, 64'h755df281d468810a, 64'h501e1140d01c3a, 64'h915df65e0},{64'h180000000, 64'h4418000000000000, 64'hf55d366b993ac, 64'h38800000c008973c, 64'h53800396000c2e, 64'he01e03c00},{64'h6001000004000000, 64'h7000000000000014, 64'h9aa9c810594b1, 64'h603017919a1e4056, 64'h5fa834f3b7a514a0, 64'h14a5e5007a},{64'h8000002000c0, 64'h3000000000000000, 64'h31959a5b663e300d, 64'h5672dceb4c297477, 64'h786380047376dc3b, 64'h638006ae1},{64'h30000, 64'h28000000001000, 64'h8bb2aba45ea00, 64'h6ae0009448e51e, 64'h15000000000eec, 64'h1a5c001180},{64'h2010030000, 64'h3000000000001014, 64'h892b002ac30b8a9, 64'hdd10d77578c785de, 64'hc84c23c72a8f178d, 64'hee445045d},{64'hc0, 64'h401b800000000000, 64'h165164db57b962b2, 64'h72c09dbd000303, 64'h5bab04000, 64'h1a580072c0},{64'h2000000000, 64'hf000000000000080, 64'h89e154939e315, 64'h2300432017000000, 64'h1d2000004e9149d, 64'h1d363d8000},{64'h800000200000, 64'hb000000000003000, 64'h119e19278e980b, 64'h5bfea63080005a, 64'h498005e7184308, 64'h1a67a20000},{64'h3000040000, 64'hb000000000001008, 64'hbdd07d124c059805, 64'h9c69fe05cf41705e, 64'h3d9daf8676000ee7, 64'heeef85074},{64'hc000000, 64'hf151800000000008, 64'h9bb5967466102, 64'hdc02f23910800442, 64'h78000000f4000559, 64'h8dc4769f7},{64'h3000000044, 64'h7000000000000010, 64'h613475a3358a180a, 64'ha2190001720005e7, 64'h7a948005ac009a5f, 64'h794},{64'h1060000000140, 64'h1000, 64'h8ed17e192c51c200, 64'h7d4fa0000e000525, 64'hc46d46168f89ee8a, 64'h1d1e3d3861},{64'h4000000, 64'h300000000000000c, 64'h7116caeb4c1421d, 64'h4b3c15bc0000043c, 64'ha91696400000024f, 64'h7250},{64'hc00000000000, 64'hf000000000000000, 64'hcb066d045621d, 64'ha9760e5d0db97000, 64'h9c0600073189cc28, 64'h21e8},{64'h300000008000040, 64'hb000000000000000, 64'h2b136565182e8f02, 64'h52f780560005e1, 64'hbdd742f680248178, 64'h8af2f15a0},{64'h8000000, 64'h420000000000000c, 64'h2c57a29ab84df872, 64'h699000ba800302, 64'hb00180030959c000, 64'h1d600752be},{64'h3000000040, 64'h3000000000000000, 64'hf884ae8f15ae00b, 64'hf452a00173000753, 64'h1ac0005e61700ce, 64'h1d0a946b00},{64'h1180020000, 64'h3000000000004000, 64'haa31d78a5f241, 64'h498c42b0c14b8693, 64'h2c3116a0c45a8c17, 64'h568b0aaa},{64'h8600000, 64'hf01a814000000000, 64'h620d9bdcc90d381a, 64'h5dda6207283506, 64'h88c48000f00c11c0, 64'h181890601},{64'h10000, 64'h840a000000003000, 64'h2f09bb2abb290f83, 64'h9169200177f49510, 64'h3c0bf13b8, 64'h91d282500},{64'h8000000, 64'h4200000000000000, 64'h2509baa4fada0374, 64'h9414125000000681, 64'hd4e6135398250e58, 64'h968003864},{64'h4000020000, 64'h8200000000003000, 64'h468b4358f74e3782, 64'ha0140430c04253c8, 64'h3dbe91b6fa03c03c, 64'h1cfc613c1d},{64'h4100050000, 64'h432882c000003000, 64'h179b58f709385d, 64'h94d2e48c5cd23000, 64'hfc940001924a1d06, 64'h19dc5818e2},{64'h0, 64'h5000000000008, 64'h31537558b7c92100, 64'hf0f44548a8c60f4, 64'h200000021e6203d1, 64'hc40006af6},{64'h400000100c0, 64'h2c00000000000000, 64'h2f0b43e75a3af194, 64'h35dc000ee6ef11d, 64'h94218796b10ab770, 64'h1d51257544},{64'h400000000080, 64'h7128000000000000, 64'h8fc9bad11555830b, 64'h3bb8fd6f35772d, 64'hddcb000479b591f8, 64'h1be8006ae8},{64'h300000000000000, 64'hc400000000000000, 64'h1385d4bab101a3, 64'ha3000001a5c31238, 64'h14a7a309200024b, 64'h8e8000160},{64'h23000000000, 64'h3107000000000008, 64'h2f4d54455c02d802, 64'ha50c2e9418922244, 64'h884b000249e93d5f, 64'h1c5800699e},{64'h30000, 64'h3015824000000008, 64'h1144eb7b0e9813, 64'hc738a6da7c0c22a, 64'he14d8cc018a6dc20, 64'h8b0003bbb},{64'h460000000000, 64'h405800000000000, 64'h166a1ec9c5d594, 64'h7a248308ee221094, 64'h11100067746e488, 64'h918000000},{64'h0, 64'h5800000000002180, 64'h47089ca9008ed8ac, 64'he43d8000f6000443, 64'h2896800694d1c969, 64'hc2ef4a5ad},{64'h10200080, 64'hf000000000000000, 64'h78d28d16f731500d, 64'h70f4a6e29e35c9, 64'h906d0007471e0690, 64'h4787},{64'h300000000400000, 64'h3000000000000000, 64'hc862f55a9e115, 64'h4fb746b7b4b000, 64'h1c94002cee8d108, 64'h16ba30140},{64'hc0, 64'h3000000000000000, 64'h878953e8e0d50204, 64'h5be12400000731, 64'h95138b345b2bc598, 64'hc2800166b},{64'hc01000040000, 64'hc400000000000000, 64'h5c529adaa821f865, 64'h4044e4e5c3f97c42, 64'hd84b00022b0bcc2f, 64'h5687b6645},{64'h20000, 64'h3017810000000000, 64'h164caf35c54313, 64'hee1cf079672c, 64'h30828cc28, 64'hb50000000},{64'h860000000040, 64'h3000000000004000, 64'hba0e7c2b3b02580a, 64'h5b4001740002eb, 64'h7d4a05f305eaf538, 64'h11c00759b},{64'h1000000000, 64'hf00000000000000c, 64'h495282d8d106980d, 64'h62164328c00a771c, 64'h5dac4b23042c97a4, 64'h1cb926743e},{64'h80, 64'h5c1880000000000c, 64'hbfd79a5165bdb2a5, 64'hfebad7b800531, 64'h24183582d58e4000, 64'h1acb005336},{64'h40, 64'h26016000000000, 64'h17a25b343e4300, 64'h4f400000000507, 64'h4524017a921240, 64'h1448003c00},{64'h40800, 64'hb000000000000000, 64'hd4f6c1121298303, 64'h25a0d40bf4997a, 64'h928001004941a8, 64'h400002512},{64'h40000c000080, 64'hb000000000000000, 64'h640b439967ce1704, 64'h397d10c4000129, 64'h9ac00399001a20, 64'h321910000},{64'h18400008000000, 64'hf000000000000000, 64'h2517a2448c0e181c, 64'h1452919c5f894246, 64'h108df50efb04c940, 64'h65284028a},{64'h400000001000, 64'h2d7a800000000000, 64'h31899ad4f8869002, 64'h22a00091e98a1e, 64'h64c409925143c4c8, 64'h6300022c2},{64'h20000100c0, 64'h6000000000000, 64'hbc0f459ab84aea00, 64'h8ac000f5, 64'h100000009a2f487c, 64'hfa0},{64'h2000003000000000, 64'hf000000000000000, 64'h18577086ac01f80a, 64'haa4fae811f87a0f4, 64'haa01000754a0d1e7, 64'h16c80524be},{64'h80100c0, 64'h316a828000000000, 64'h19d3662577b9311a, 64'h72dd09abc675bd, 64'hc0568002d4001a10, 64'hd05},{64'h1000000c0, 64'hf000000000001000, 64'ha48e62ef5506180c, 64'h24f1674dab800249, 64'h17cd61d1d, 64'h1a6c000000},{64'h40, 64'hf000000000003008, 64'h1514bbc2ec02581c, 64'hcc74be1dce0cc245, 64'h4c2f0001980014d8, 64'hef6906a11},{64'h500000000020100, 64'hf018000000000000, 64'hd011756931b1784d, 64'h303ba47c06498171, 64'h2ac0001ccec920, 64'h8b4007040},{64'h300800000000100, 64'hb000000000000000, 64'h134f8de550c26053, 64'hc60184a40604d01d, 64'h39115155e94b4878, 64'h8e8003ca1},{64'h400000001800, 64'hb14909e000000000, 64'h13462116deab02, 64'h5b2134f6529b96, 64'h51188006958c56c8, 64'hf200038c2},{64'h0, 64'hf014000000002180, 64'ha5da139099813, 64'h698e586d5e33d8, 64'hac1a16b3d8e58950, 64'h11edd2efe5},{64'h10030040, 64'h6c00000000005000, 64'h5dcb835ea9c98275, 64'h14100116d772df, 64'h2a8007472cd108, 64'hf2e9752e0},{64'h400860000000000, 64'h3017800000000000, 64'h962855c0af81c, 64'hd33a60019a00044c, 64'h63c0030b89f0b9, 64'h5cb0},{64'h6000000008000000, 64'h3000000000000004, 64'hbf1680071c0e5815, 64'hd3681ceda4915692, 64'h868d80018e0d59d9, 64'hef0002ed7},{64'h300000010000040, 64'hec00000000000008, 64'hbd888e2ae641f3a5, 64'h665ddbfd732ff72d, 64'h54bb4005bcbd0c2c, 64'h16780075da},{64'hc0, 64'h400000000000000, 64'h4a53bd5710b9007d, 64'h5ca308940005e9, 64'hd8000002ea000590, 64'hb00001965},{64'hc04000000000, 64'h3028000000000004, 64'he42e93b815891, 64'h425fe00144b586b0, 64'h305e8c24f, 64'h936f772fc},{64'h400000000050080, 64'h7000000000000080, 64'h90158d9e4c492ba1, 64'h49043c30d0f473, 64'h1d167d1960011f8, 64'h180759c900},{64'h41000000c0000c0, 64'h7000000000000004, 64'ha0d375417c2a120b, 64'h4975fb7c1a862251, 64'h957c5e1dc8a25244, 64'h167ae0513b},{64'h20000030000, 64'h2a000000000000, 64'h138a5c85deaf00, 64'h6840009ac00000, 64'h2c00000101497a10, 64'h1458006a0a},{64'h1000000000, 64'hf000000000000000, 64'h28ca80828c2a430a, 64'h4e1944a16f8a35be, 64'h400001802014ac, 64'hc8d241480},{64'h11000000c0, 64'ha6f6000000000000, 64'h7457aaa91b0e4913, 64'h28c621ac8ab8f247, 64'h7463a321327300a5, 64'h4ab9d509e},{64'h0, 64'h417000000000000, 64'h1fd29b5e8ba6aba3, 64'h953082a80000021f, 64'h580000024a2f8c28, 64'h1110944442},{64'hc000040, 64'hc400000000000000, 64'h114ad1754a7073, 64'h14757a0800000479, 64'h139b415e3050bb0, 64'ha0000000},{64'h300004100000000, 64'h3000000000000014, 64'h1ecf4466c0c0b869, 64'haac5a2b5d04ae674, 64'ha16ff032decd817f, 64'h3416015b8},{64'h200003000000000, 64'h4014000000000000, 64'ha8d59e1edb2ef272, 64'hcc39877cef084132, 64'h1a6f8c000001a6d, 64'h1520005360},{64'h3000020000, 64'h7000000000000004, 64'ha254ace3695d4813, 64'h53198001d2f97018, 64'h402a8006b1178ef4, 64'h247a},{64'h10000040, 64'h3009000000000000, 64'h30d5b61f112d83b9, 64'hc564000000739, 64'h4599000682001a00, 64'hc40002466},{64'h501060000000000, 64'h3000000000000004, 64'h61cab8a0c04d0b71, 64'h16320458b81902e0, 64'h14c4cd0061e0a8a1, 64'h270b33bd4},{64'h300000000000000, 64'hc224000000000000, 64'h116ce89b4af582, 64'h5dc000dd800478, 64'h2cf6e2f45ed60000, 64'h1ac8002557},{64'h4000000, 64'h8600000000000000, 64'hf92174059a2b3, 64'h815b300040000268, 64'h114000450001cb3, 64'h959352580},{64'hc0, 64'h3000000000000008, 64'h364ca3aca4c22102, 64'haa754014000003d9, 64'hb5f353a4cd41a3, 64'h6d0d169b0},{64'h4030104, 64'h3000000000000000, 64'h61719c9b07dd2871, 64'h3530b75513c00129, 64'hf09c638c000eaa, 64'h4c80052f0},{64'h1000000000000, 64'h3000000000003000, 64'h274d439900b26289, 64'hec44f78cbd000306, 64'he8000003117b0ea9, 64'h1a0d833bc5},{64'h1000000080000c0, 64'h0, 64'hbbd137b3e7154, 64'hf767700000000693, 64'h8dc005a20016f2, 64'h176a2e0000},{64'h460010a, 64'h3000000000000000, 64'h8ff070811c20b849, 64'h5852bbd37fc580f5, 64'hd88db3c2c4160ba8, 64'h8d90f678b},{64'h21840, 64'h8000000000000000, 64'hd2517d54b6a12c83, 64'hff2ec000936e5a53, 64'h1c019cd694e91d1a, 64'h1d30ae39a6},{64'h6000000000000000, 64'h5c18000000000008, 64'h8fd24e14b6bd88bc, 64'hd6e2da40006b1, 64'h2b243ad476eb51d0, 64'h601a},{64'h3010000000, 64'h3000000000001000, 64'hcd50939b37b2e2a1, 64'he4537a2087f7d01e, 64'h139af55a2df544e, 64'h124f360000},{64'h0, 64'h8200000000000000, 64'h176a5f6acd828b, 64'h52a00000000000, 64'h940000068e000000, 64'h17068d51ae},{64'h5000040000, 64'h3000000000000000, 64'h30d24864a181c259, 64'h75ed380674d252, 64'h1488206a100096c, 64'h5200009e0},{64'hc000040, 64'h3004000000002010, 64'h45556ce57b055861, 64'h251735188005bf, 64'h343634d32a331a20, 64'h924003c9d},{64'h0, 64'hc600000000000008, 64'h864b8366e0d180bb, 64'h44e4940000012a, 64'h1d5001752300928, 64'hbe22773b0},{64'h4100030000, 64'h300b000000000004, 64'h107cdcd626f241, 64'h85cea05092e825e4, 64'h3c00000072e7459d, 64'h1793984450},{64'hc000080, 64'h130000000000000, 64'h2b895bd0eb564100, 64'h6f683001953912ed, 64'h2c4e5c0a5, 64'h5700e6740},{64'h8000000, 64'h0, 64'h154be2e1aa81ba, 64'h45b2294d88a3bc, 64'h10a4bc000, 64'h9788b25e0},{64'h40000c0, 64'h3000000000002000, 64'he70a43eb34d9c015, 64'h7e3990011e80074b, 64'h1c50551a89f82f2, 64'h1524d41a80},{64'h200000010000000, 64'h4200000000003000, 64'h620a4b9f48dd8083, 64'h98165001cb80c320, 64'h1484005c0a69703, 64'h1455241960},{64'h3000000040, 64'hc400000000000000, 64'h7194ac5cf82540b5, 64'h90000008a0d0681, 64'hc300053c001a0d, 64'h14f1c753c0},{64'h20040, 64'h7000000000000000, 64'h8b0a43aec4d22305, 64'h22d8b4c87462e1, 64'hd0e58000000010b8, 64'h37c8},{64'h100, 64'h3000000000000008, 64'hd01784d8a08963a9, 64'h3680cd09600006b, 64'hc800032e99d30, 64'h1acc1247b0},{64'h63008000000, 64'h3000000000001000, 64'h8e4c4b9f184a770d, 64'h72d345d52f95f2, 64'h32314515afd7c, 64'h9ae3a5f40},{64'h1023000000000, 64'hf000000000002000, 64'h78976a6d55019414, 64'ha075526560800450, 64'h19d72c6101cd6e97, 64'h6d62975cb},{64'h24008600000, 64'hf000000000000000, 64'hba355165ae904, 64'h9e3c38d693125186, 64'hbd1e438d7864cc, 64'h3060},{64'h300002000000000, 64'h7000000000000000, 64'h1e95b51510b22013, 64'h845bce580000072c, 64'h44ef4005a61f0f67, 64'hc87d0320},{64'hc00000010000, 64'h8000000000000008, 64'hfba50b54e3693, 64'h2eabd980495128, 64'h6d4780045d590000, 64'h4b0005db4},{64'h100000000000000, 64'h3025800000000010, 64'ha615b224f1867861, 64'hb30e7982c6983cc, 64'h19e74a724e44f30, 64'h1468000d10},{64'h100000000000000, 64'hb036800000002000, 64'h1545df174e160c, 64'h474888bb622000, 64'he6c6c490900000, 64'h1d35e223e0},{64'h4000000400c0, 64'h3000000000000000, 64'h49d34d64d039e251, 64'h5c89d466688691, 64'h9380075bb4c8e8, 64'h5c0b723c0},{64'h10000, 64'hc400000000000000, 64'hba9042989bc9e3ac, 64'had5088f9bee8451e, 64'h1c600075a001a83, 64'h19b4000000},{64'h300000000000000, 64'h3028000000000010, 64'hb90e64653a82c1b9, 64'h2500014aef5180, 64'h1d2c31060000188, 64'h16cb3609d0},{64'hc00000000000, 64'h400000000000000, 64'h9ae1ae84ac1ba, 64'h69d1b0dd8cc462, 64'h2063800523320000, 64'h8b0003a23},{64'h0, 64'h4600000000000000, 64'h4b63d540da6245, 64'h850b06142c179436, 64'h1a6c00312001d49, 64'hc880044e0},{64'h0, 64'hc34900000000000c, 64'h18c8762359aac285, 64'h24b9dd74061504, 64'hc8318005e2001788, 64'h1d0002f9b},{64'h0, 64'h200000000000000, 64'h80ea4195bda625a, 64'h2ded39d600069a, 64'hb19d00073b590038, 64'h5780065ae},{64'h0, 64'hc234000000000000, 64'he94b852d79b14293, 64'h738e1042b8c114, 64'h9790f72fe748d8, 64'hef91b74c0},{64'h0, 64'h41b018000003000, 64'h96c2f554a6f45, 64'h72ce10bc800754, 64'h11f0d472e608c10, 64'h152fab71a0},{64'h110c000000, 64'h3006800000000000, 64'ha696525f484a6e0b, 64'h9d8bdeacc800001c, 64'h3100013f7, 64'h1cc0000000},{64'h1010400000, 64'h3000000000000000, 64'hbe08b0037c51c399, 64'hc8747492c300018e, 64'h14f30018cc01704, 64'he0160380},{64'h200000000030000, 64'h3006000000001000, 64'h84aace8b6ef0d, 64'h490c41288b463432, 64'h8ae3d396128318, 64'he3e2d3800},{64'hc0, 64'h8026800000000000, 64'h4510955f19b9414d, 64'ha0024431a000068d, 64'h8a800756001d5b, 64'h80},{64'h1000000000, 64'hb02a000000003000, 64'he8ce8c2f36055804, 64'ha41502b924000490, 64'h57801033905d37, 64'h9b6fa15a0},{64'h20000, 64'h3014800000000190, 64'h176c66a651f691, 64'h9d396369d55c5000, 64'h4d6139d3c60006d3, 64'h11d4db9493},{64'h8000000000000, 64'h3116800000002000, 64'h105cc4ec4aa303, 64'h24a000f01d4180, 64'h1637ae800000000, 64'h114c003ba0},{64'h3000020040, 64'h3000000000000010, 64'h6252b0284c2898a9, 64'hd63ca000bd6de307, 64'hb4c8800322be0f6e, 64'hf6b0012d7},{64'h10000080, 64'h4600000000000004, 64'h25497e1125b2eeac, 64'h2f0290c4baae972d, 64'ha52100007291cb38, 64'h3ec31033b},{64'h860000000000, 64'h20b800000000000, 64'h838f6616eaa633a4, 64'ha4090a90f304a016, 64'h7505800679a3fc8a, 64'h107800094a},{64'hc00000000000, 64'h822a000000000000, 64'h485762152ac57385, 64'h480d84891d240531, 64'h39b2e4f12, 64'h0},{64'h300000000000000, 64'h4400000000000000, 64'hd1177ce92082188d, 64'h454ee2dd116e4510, 64'h8fc2024e0016b3, 64'h0},{64'h0, 64'hc200000000000000, 64'h75576c6d21d60274, 64'hd6684359ac08452a, 64'hfc000006b2498931, 64'h23d8},{64'h300000000010000, 64'hf02b000000000000, 64'h2797ac69273e700a, 64'h3523e4d542529306, 64'h4575d83062079d6d, 64'h172b5125cd},{64'h0, 64'h84170d0000000000, 64'h91497ae2a9b6f6ac, 64'h75a90cbd3ad13c, 64'h1d7cc83a25e8000, 64'h1c724666d7},{64'h200000000000000, 64'hc20680000000000c, 64'h8b579a5f6a491572, 64'h4420008e800170, 64'h791962751a8b4290, 64'h10fa8e22d4},{64'h300000004000000, 64'h400000000000000, 64'h89cf95e965ba096a, 64'h30b18d3d0005c8, 64'h9dd56f2074b94c8c, 64'h141a1c5b28},{64'h0, 64'h8619800000000000, 64'h1653d69ba2826b, 64'h67000000b787c000, 64'h10bac67402178d, 64'h1a707d65e0},{64'h0, 64'hc09a800000000000, 64'h1488dca121816b, 64'h6d10c001ce387000, 64'hefa32000001d00, 64'h1d30004640},{64'h0, 64'h200000000000000, 64'ha8b5921d2a244, 64'h71aea5cb387000, 64'h9d50026780008dc, 64'h682c},{64'h40000100c000000, 64'hb00000000000000c, 64'ha08e5aa6d652a204, 64'haf4fda0d3b970020, 64'hcc8df982e04dcc17, 64'h1d5d717632},{64'h1000004030000, 64'h8000000000000008, 64'hb0155a62f75e936d, 64'hfd5c1059d5f8c58a, 64'hec643ae695bf5d6a, 64'h163000323b},{64'h6300800000000000, 64'hf016000000000000, 64'h7a56ba1eb8c2ad04, 64'h4a0c6a253b9e9510, 64'h1fd85c3601798e58, 64'h397},{64'hc000000, 64'h18824000000000, 64'h16a4eafbc1a200, 64'h45bb79d5006000, 64'h4c0000039ab7d698, 64'h8a90f3a46},{64'h10000080, 64'h4000000000003000, 64'h4e5aa707a121a5, 64'h886a15d4c8000751, 64'h4dd80002ec000b21, 64'hd7a43986},{64'h100000000030080, 64'hc000000000000000, 64'h86d48e18b54e0e4d, 64'h4545abe4545cb491, 64'hf457c454d40e9350, 64'h17ea6645ab},{64'h6000000000000000, 64'he42a800000000004, 64'h904d7c5c98226b55, 64'h1b500090800490, 64'h1f4985d0b0000000, 64'h149a49453b},{64'h40080, 64'h300000000000100c, 64'h16ba414c21cc69, 64'h748ae7c2c526bbb, 64'h9d00af600be5228, 64'hf0caf3ab9},{64'h6000800000000000, 64'hd4800000000004, 64'h5a538b20b939e000, 64'h484000000002ea, 64'h7f748003230c5238, 64'h1d1853dbb},{64'h0, 64'h3027800000000010, 64'hb616b8d880c24049, 64'h32000001c880d5bc, 64'h7c99000000000251, 64'h979da15fb},{64'h1400008000000, 64'h7018000000004000, 64'h16bae951b11149, 64'hdc549a848b2a1000, 64'h98bf1ed25fa7c8d8, 64'h45e0fbda7},{64'h1020000600080, 64'h3000000000000000, 64'he58a5b69184df561, 64'h972459233d000445, 64'h9d7b8a1a98ee93b, 64'h1448b8676c},{64'h0, 64'h4600000000000008, 64'h88976c58b5228182, 64'h548a75520006b0, 64'h68e215a2c, 64'heb3495cb0},{64'h12e20000000c0, 64'h3000000000000000, 64'h7929d2ce0a1e049, 64'h832446284f8b9509, 64'h53dec2935, 64'h9118e31c0},{64'h10000040000c0, 64'hf000000000000000, 64'heb099a9159468205, 64'h7a26b02800000253, 64'h18e1a4447b27ce89, 64'h1d68006a39},{64'h20100, 64'h5600000000000000, 64'h7b979a20c1c5e103, 64'h1d6ef9681, 64'ha57e80044e885468, 64'h1236fd0a68},{64'h2000000000000000, 64'h5800000000000010, 64'h7b8e78e0a12ee04d, 64'h26a4b89aa0b074, 64'h7a000005e4ec0000, 64'h1078005f54},{64'h44000000000, 64'hc200000000000000, 64'h5a48ae253a3ac37d, 64'h3a1b434c108da2de, 64'h1990005cba0fcef, 64'h69c0},{64'h30000, 64'h400000000000000, 64'h129d62c0dae055, 64'h875c0001d6400738, 64'h1d30005caa98ef8, 64'h1d280c7140},{64'h0, 64'h580000000000000c, 64'h127ba110d94242, 64'hf01d4752, 64'hd1972f680000000, 64'h74d0},{64'h800000000000, 64'h300000000000400c, 64'h16585cd05098a9, 64'hb34945bc0e0002e0, 64'hc40000072fe60b20, 64'h4b400757e},{64'h100, 64'h4000000000000000, 64'hfa0d7214e01b4, 64'h5fa0017d8003cd, 64'hf40bba2506000000, 64'h5069},{64'h218001000000000, 64'h7000000000000000, 64'hb60a5b83490d9813, 64'h91396714000005c8, 64'h1d741cb226297ed, 64'h1635e75ca0},{64'h40, 64'h7000000000000000, 64'h80e7c6d754a620a, 64'h45513b596f0003d3, 64'he00003a28ec36b, 64'h11db4522a0},{64'h3000000000, 64'h25000000004000, 64'h9bc5107d26173, 64'h2ce000bab4f000, 64'h11c0396001d5c, 64'h14b4007480},{64'h500004000000000, 64'h3000000000000000, 64'ha60e92139a1a9, 64'h66000000c8c00240, 64'h172e2d08a00018e, 64'h10f8000780},{64'h1001000000000, 64'h3000000000000008, 64'hdd8d40c31c3940b1, 64'h725129282c3ac508, 64'h4c00000191eb1357, 64'h4b775fba},{64'hc00000000000, 64'h400000000000080, 64'h178a6d393d155d, 64'h52800121000000, 64'h14c28c0bb000000, 64'h124d278000},{64'h2004000100, 64'h3000000000000000, 64'h8e01a6184c489869, 64'h3c48b028000000c7, 64'h1d04005d20e9806, 64'hbb3a774e0},{64'h8000000, 64'h300400000000400c, 64'he5899a9cf0c498b9, 64'h1548f4248a077722, 64'h283600072e1dc079, 64'h3eedf30be},{64'h2000000000, 64'h20480000000000c, 64'ha74f656938dd6eb4, 64'h8e264000993ad542, 64'h6d508005424c0997, 64'h1500003b54},{64'hc00000020000, 64'h2c15800000000000, 64'h5e558e197749f412, 64'h8524e00150c0030a, 64'hf4f6f2f2fdce85c1, 64'h5129},{64'h0, 64'h4200000000000000, 64'h11bd94b14a037b, 64'h2300000042800000, 64'h94800694001cbd, 64'h1ac8003ac0},{64'h4000000000, 64'h300000000000000c, 64'h8705541309889, 64'h140a5152583000, 64'h910bb000000644, 64'h17a0006930},{64'h300000010050000, 64'h3000000000000000, 64'hc8559098d0ccb841, 64'h955e831c9f488, 64'h2dace460000018e8, 64'h19100031d0},{64'h40, 64'h9a0000000000000c, 64'h34d782275101781d, 64'h2d51a0680d0003a3, 64'h446bba71aee9c29a, 64'h1d6c1648d0},{64'h300000000000000, 64'h228800000000000, 64'h134d1ab7b2ee94, 64'h8e44f88400000000, 64'hf17ec3b44e639791, 64'h7e0f73183},{64'h10000, 64'hc600000000004000, 64'h30484adea8c1a274, 64'h674cd09acb925c, 64'h5a713226400107c, 64'he65700443},{64'h0, 64'h8624800000000000, 64'hbaddb674a6162, 64'h9744e0006d400018, 64'h95c839730200113b, 64'h17298573ae},{64'h400000004000000, 64'h312845a040000000, 64'ha609761a49871, 64'h3bfd01a7800668, 64'h3057c00000000000, 64'h2000754d},{64'h10000080, 64'h3000000000003000, 64'h5bca402760d09859, 64'h63000000003c1, 64'hc000004fabc0000, 64'heaef42d4a},{64'h40000, 64'h3000000000003000, 64'h79d75096e0a49879, 64'h773a2714256fd3a2, 64'h1419ea5f8dddcc7, 64'hb8f763d40},{64'h803004000000, 64'haa06000000000000, 64'hba0f4c5576ca760b, 64'h5fb7a8e5af173e, 64'he1d01fd039bc5d74, 64'h1728093fa7},{64'h0, 64'h398a8140000000, 64'hb78fbd54b6d92c00, 64'h3a20000000038a, 64'h651d8210dc000c8c, 64'h68ab},{64'h0, 64'hc400000000000000, 64'h5d4c7054d04ac3ba, 64'h396ea00000038a, 64'ha9c6000748001d40, 64'h65},{64'hc0, 64'hc200000000000000, 64'h3a9064dca04ac2ba, 64'h4d24cd10750e569f, 64'h340000045a884933, 64'h1aed},{64'h402000000000, 64'hc00000000000000c, 64'hb9c695bc15273, 64'hac01283907000000, 64'h25050004d79f422f, 64'h1b9800243a},{64'h300000000000000, 64'h3000000000000000, 64'h6c936523212de102, 64'hae3aa0c5a1800472, 64'h149e3a48c8c4ef1, 64'h1bbdb33bc0},{64'h80100c000000, 64'h5207000000000000, 64'h5e549e152859edbc, 64'he9519000c1298074, 64'h352480052b6094c6, 64'h124a48532a},{64'hc020000, 64'h8200000000000000, 64'had084b1f7a556a8d, 64'hb04731b11e50c228, 64'h5c0000071e0003ba, 64'h15a80074fe},{64'hc00000000000, 64'hc000000000000000, 64'h178a16e15aa184, 64'h54000000000264, 64'h1c88007250014f0, 64'h98aa20000},{64'h400000020006, 64'h3000000000000000, 64'ha8624580cc0e490c, 64'h2f30a5f09955275b, 64'hd544957543e499a8, 64'h1c90102aec},{64'h80, 64'hc01600000000000c, 64'h35cb8c1556a12f94, 64'h3c29f46b86124f, 64'h64eb0863c2760000, 64'h6b27e677d},{64'h300002000000000, 64'h4205800000000000, 64'hcd13aa5cf9511763, 64'hfd674001b2000176, 64'h98927662447f494d, 64'hfc800676d},{64'h200000000000000, 64'h820000000000000c, 64'hd40ba35e88caea75, 64'h6ecdc5a8376307, 64'hdd4af7748a075b98, 64'h5e9d},{64'h418800000010000, 64'hb000000000000000, 64'h6947de53aae0d1b, 64'h2c000bd41151a, 64'h8ae46f5d1506a0, 64'h1914000000},{64'h440000000000, 64'h7000000000000000, 64'h545678c12b8a180d, 64'h275e40000d43b2ac, 64'h953500074f35e7ba, 64'hab8004d49},{64'h1000000000, 64'h3038800000000000, 64'h2e0a5b2d744aa204, 64'h2f0440019d12724e, 64'h5d80069c304c75, 64'h1f90},{64'h400000000000, 64'h702a000000000000, 64'hb995bd9d21bd800c, 64'h31c398c60005e8, 64'hadd139d265bd0c70, 64'h7580074c3},{64'h200000000000000, 64'h20680000000000c, 64'h5150a49f7b226b53, 64'hb328a501a01451ee, 64'hc2cfc1f86cca09, 64'ha31b23050},{64'hc0, 64'h621a000000002010, 64'h7b0db3a53ade087a, 64'hec3646b4d9000699, 64'h91d5683342670d09, 64'h1a85702ed7},{64'h6200000000000000, 64'h16812000000010, 64'h115ddcf84a7400, 64'h766ca000e8b655f8, 64'hc77a7613d4000f43, 64'h5bfb},{64'h100004000030000, 64'hb02a000000000000, 64'h126d430702381d, 64'h778127e17ee54000, 64'hf56590260008df, 64'h1d00154b20},{64'h100000000000000, 64'hf000000000000000, 64'ha889761556a2420c, 64'hfc544a6d78dd13fa, 64'h88fef2268a0018f1, 64'h16f9fe044c},{64'h0, 64'h82340aa000000000, 64'h129dd706da2972, 64'heb5d63ace5af1620, 64'had86b91477001788, 64'hbb3111d4e},{64'h1000000000, 64'h12340a8000000000, 64'hea0b6e212ac553b3, 64'h2d7510007e0001f8, 64'h2da68e668e3edd26, 64'h74e0},{64'h8000040, 64'h7038800000000000, 64'h9a8a5de8fb31c00b, 64'hc624deb187ac21d5, 64'h144b1158c00134a, 64'h526b6220},{64'h106, 64'h226000000000000, 64'hddeaa36f04bab19a, 64'h2ae0010755745b, 64'hef1563b0000000, 64'h11d1af4680},{64'h0, 64'h7000000000003000, 64'ha3d26d50a131c11a, 64'h465d25f000000530, 64'h241d80028c000c11, 64'hd9d456899},{64'h0, 64'hc205800000000010, 64'he4c64c1dae284, 64'h591f84b12a8001f0, 64'h87b974b24d47e2, 64'h8a9352e10},{64'h1805010030000, 64'h416800000000000, 64'h99be1693a9143, 64'hed44f4c43bdcc128, 64'h88f69ec5cb731cbd, 64'h15ad33542a},{64'h0, 64'hb035800000001100, 64'h70c6c5f6a826912, 64'h68044c2800265, 64'h659a9530000000c8, 64'h1d76a2f240},{64'h100000000000000, 64'h703a000000000000, 64'hb9c157132400b, 64'h10c3593ea0d0cc, 64'habe0f3ac000f08, 64'h6c00041e0},{64'h1000000000080, 64'hd018000000000000, 64'hb7caab5d21d2c014, 64'h58c0019d2c61af, 64'h905e2c55077ac910, 64'h17004f3d67},{64'h100000010a, 64'h62a000000000018, 64'h72ea5bee9449b583, 64'h9a4b27312caff3d5, 64'h1b365848cbdcfec, 64'he90005cbc},{64'h200000000010000, 64'h37000000000000, 64'hc2d38a2af5c9b400, 64'h10622001bb73b6a1, 64'h19bbc176760c0e33, 64'hd8941b07},{64'h46, 64'h5025000000000000, 64'he9f1bc9cfaad300b, 64'hd11ce00179000035, 64'hccd98eb1d6368d78, 64'h1474da0786},{64'h18000000000000, 64'h8400000000001000, 64'hb5898bd706364ea2, 64'hc1750001d438c176, 64'h39354fddae001a70, 64'habc232661},{64'h0, 64'h8435000000000000, 64'h175ba55a41218d, 64'h425e8bacc700024f, 64'h195a94631a001589, 64'h56a5},{64'h300000010000000, 64'ha800000000000008, 64'ha8ca831716ca6103, 64'hf48d63a0000021e, 64'h5d369b18ca90d91, 64'h1d75},{64'h3000010000, 64'hf000000000002000, 64'h1e9175aed78e180a, 64'h3d8790a2d6a442, 64'hb4c4a221f95a8d9c, 64'ha35913222},{64'h1000020000, 64'hc000000000000000, 64'ha0c9629ebadaed94, 64'hea0c4120d96d95fa, 64'h1bba845b2000d0d, 64'h1ba0003d20},{64'h400000000000, 64'ha23b000000000000, 64'h17935d3ab1020a, 64'hf94ca001b2f766ee, 64'hc9350003d59acfe9, 64'h5000740d},{64'h101000000000000, 64'h4600000000000000, 64'h74c93eabb290284, 64'h996cc70db2b616a0, 64'h112cf595131ed140, 64'h11400002b7},{64'h101003000000000, 64'he000000000002000, 64'h138ae9595aed43, 64'h801d4bc586a27545, 64'h89914006b3b05a2c, 64'hff6c658e8},{64'h8000000, 64'hb019800000003000, 64'h97a971a8e9814, 64'h1d7e8d910001f6, 64'h9dd5f2269a000000, 64'h188f1f1d63},{64'h2, 64'hf027000000000000, 64'h3f2d4d14b186d804, 64'h41e63d0720a751, 64'h1619fe31e620000, 64'hff1fd0000},{64'h2000030000, 64'h3000000000001000, 64'h5c0e7cd096d2b213, 64'ha13442cdd65b2338, 64'he988d763bc0e9635, 64'h135ee735c8},{64'h100, 64'h8627056000000000, 64'h24097e23695e6daa, 64'h90304498abcd944f, 64'h12ca5510a000a28, 64'h14c9274b40},{64'h10100, 64'h3039090000000000, 64'had5175d8d54ea904, 64'h2d00000174e2d675, 64'h9aa56450204a35, 64'h15aab122a0},{64'h1002004000000, 64'h7035000000000000, 64'h84ddcfab22013, 64'h661f9730ab956000, 64'h89b336573b2692cf, 64'hac000264a},{64'h0, 64'hb035800000002010, 64'h4914aa18d8cde112, 64'h1224800090800252, 64'ha80000066a064f6c, 64'h99c356834},{64'h1420010000000, 64'h400000000000000c, 64'h16a2e54bb9227c, 64'h90507000c88004fa, 64'h5c33a6b2e1e4ac89, 64'h135a6a2b13},{64'h1000000100, 64'hf000000000003000, 64'h4cc84b611a59821a, 64'h2d5fc5f89997e3a3, 64'h107deb5fcbdceb5, 64'h6c5e50000},{64'hc020000, 64'h4000000000001000, 64'hbdd38d691bb9f26a, 64'ha7245045635d15fe, 64'h107a0e2a4e9d07b, 64'h1705572b00},{64'h1000000020000, 64'hc20a800000000014, 64'hc88f9c58d825cab5, 64'h6760012cc1706a, 64'h64e30005bfc44000, 64'h19131e3a52},{64'h1000000000000, 64'h7007800000003014, 64'h5c84dd8b14ac11d, 64'hff5b200180011030, 64'h696f84e2ed001802, 64'hdcd23993},{64'h1008000100000c0, 64'h4000000000000000, 64'h17ada11a49ac5a, 64'h45b3046d0d95e5, 64'hcd9cbc1d7cd4618, 64'h6db3b06a3},{64'h10410000, 64'h4600000000000000, 64'h5bcb6c29543d499b, 64'h513d3bd46f431a, 64'h38341705af161448, 64'hb5000508a},{64'h8000000030000, 64'hb02a800000000000, 64'h8fcb7e14c85d0d1d, 64'hed53643cc750f48c, 64'h15ad46a2a7b4659, 64'h1520cc48e0},{64'h4000000000200c0, 64'h117800000000000, 64'h5fd6baaa9722419c, 64'h2d42c8d9dec28d, 64'h124cfd1f83e0000, 64'hf29801480},{64'h201000000000000, 64'hc200000000000000, 64'h17525cf6d50394, 64'h3d2ddc26867198, 64'h11140072f46d6c8, 64'h1421163230},{64'h1003000000000, 64'hb029800000000000, 64'h9b3e140a2a01c, 64'hd16ee361d5b9e1b0, 64'had113ab545000f54, 64'h1110803fc9},{64'h200000000000100, 64'h35064058000000, 64'h518dad271b212c00, 64'h74e36c3dba730b, 64'h65d04176cc3486d8, 64'ha3142450d},{64'h10000000, 64'h62585c000000000, 64'h107ce4daa13755, 64'ha63c3e989a93458c, 64'ha188b101d600113b, 64'h9b0043893},{64'h0, 64'h441802c000000010, 64'h114ce954396363, 64'h371f8c89d40eb0e2, 64'hdd127d1f28dd41a, 64'h677a},{64'h4000000000, 64'h61a826000000000, 64'hfb456d849c2a3, 64'h8f676051632c5000, 64'h54c481541e001235, 64'h1a08363fc0},{64'h1000000000000, 64'h27054000000000, 64'h40b9b649452a38b, 64'h366df4d9ba26fa, 64'hd98021b1689d10, 64'hbb1b00000},{64'h0, 64'h39090178000000, 64'h96506d677b313400, 64'h12000042ab524c, 64'ha32b52644bc990, 64'ha1ab25cf0},{64'h1000000000000, 64'h2b06e000000000, 64'he7c1a9ab10395, 64'h56a0012ca58000, 64'hf4c5afa267df5168, 64'h1bf01031cb},{64'h800000000000, 64'h4618024000000000, 64'h308a6616dc3d28a5, 64'hb3030051522a32ae, 64'ha0b40c326bd980c0, 64'h1528b82665},{64'h20000, 64'h503505e0b0000000, 64'h79909c97165d2da5, 64'h91000000e65243d2, 64'ha0108000589ed3da, 64'h951ea0581},{64'h2180000000, 64'h1c1a810000000000, 64'h7591be2d74bd7053, 64'h19b22000549d613c, 64'had51800546a799ac, 64'h5508b1b09},{64'h0, 64'h35064058004100, 64'hc7baa9bd2c800, 64'hd748a90922800000, 64'he97c2fd1ae3517f0, 64'h17f67edfab},{64'hc00000000040, 64'h400000000000000, 64'h55ce7c54b6ca7483, 64'h314f6000bf79e267, 64'h317c0673d783dd70, 64'h1803ae4f6d},{64'h0, 64'h62b85e000000000, 64'h798b8e14d926b043, 64'h99644000f58113d6, 64'hd91b00038c001d3c, 64'hd1e50328},{64'h41000, 64'h420900000000000c, 64'h4814bd95542d2c74, 64'h24c0178f3b81c, 64'h6d3821a4e08640, 64'hc2df0370},{64'h4000000000, 64'h8024866000000000, 64'h59d7861b67b1c344, 64'h1c1640019d0171b4, 64'h90578000385a1a6c, 64'hbd9792f62},{64'hc0, 64'h9e2a06c000000000, 64'h6389661d58a16abc, 64'h3468e0002c347183, 64'h1472894681b861e, 64'hb80230000},{64'h500004000000000, 64'h3b890168000000, 64'h87d24d5cf8b28000, 64'h9c00000087a40196, 64'h11d6a443e200ef6, 64'h12380022a0},{64'h40000, 64'h4015000000000014, 64'hd4e7de961b62245, 64'h694000c174a664, 64'he86cba81b2350130, 64'h7eb33533b},{64'h4000030080, 64'h2a14000000000000, 64'h5f0d5e18f75ae994, 64'h3d4280b54633d9, 64'ha09a2982684bc8ac, 64'hc057d5081},{64'h400000000010000, 64'hc439000000000000, 64'hdae18f75e6952, 64'h7f6fe0016cc0001c, 64'h8d517a2237201d5b, 64'h1d180a444e},{64'h40, 64'h4000000000000000, 64'hbad1b49095a9e283, 64'h28cb656c8cc1b1, 64'hf04090d450434000, 64'h17600009c0},{64'h10000, 64'h629000000000000, 64'hbb8dabeeb44d5473, 64'h531b70fdd3ceb26a, 64'hc4a8b622768ed0, 64'h177aea5d40},{64'h0, 64'hd4370aa1b0000000, 64'h5cd8e1ec85e684c, 64'hf774d045d381774e, 64'h6d41af869246da4a, 64'h7eba87524},{64'h0, 64'h54f5890160004180, 64'h1c54ad9cd85e784c, 64'h32464129a000c58c, 64'h1c4000710bc11be, 64'he97a98000},{64'h10600000, 64'h2b068000000000, 64'h70cf9e195746f200, 64'h62363fbe81c016, 64'had29134321c40, 64'h1c41c40000},{64'h1000, 64'h4200000000000000, 64'hd7e11685dc9a5, 64'hd28cad5d15b3996, 64'h150800466201509, 64'h14f10d0000},{64'hc0, 64'h29066000000000, 64'h70e7e188826d100, 64'h23664001be8b9121, 64'h8f000190000995, 64'h8f0356660},{64'h2000000000000100, 64'hc400000000003000, 64'ha911761156492aa5, 64'h875da761769d85e9, 64'hfa1d8000860014e0, 64'h12d40031fb},{64'h110004000000000, 64'h3b800000000000, 64'he10e66250a4e3500, 64'h7031129d200d748, 64'h74b44c3800000f6c, 64'h17409670a7},{64'hc02000000000, 64'h5400000000001000, 64'h6c89e169c5236bd, 64'h125232800d98a152, 64'hc70000596053dc, 64'hf558e15e0},{64'h40040, 64'hc400000000000000, 64'hd14f56291ba6acb4, 64'h30000001bbf453ad, 64'h160005470b0132, 64'h1187d0000},{64'h1010c000c020140, 64'h0, 64'h96514e2b0bb10f00, 64'h8f5fd87d22e1f6ef, 64'h17ec813fd9ae6bc, 64'h12d08b0000},{64'h400002014200000, 64'h8b80000000000c, 64'hbf514e26da800000, 64'h6cd9efa658a31e, 64'hf9acc00000001d74, 64'h601b},{64'h200003000040000, 64'hbb800000001014, 64'ha456ae0000000000, 64'hae74600113e403d7, 64'h11b40075c000e37, 64'hd69258f0},{64'h4400000500c0, 64'h4000, 64'h6397aa5d28800000, 64'h6d1141d5915db031, 64'hbc90c0070536aed8, 64'h7657931e2},{64'h500061010000000, 64'hab800000000008, 64'h2e095e271c425500, 64'h9941f75c0c017030, 64'hff4002f35a20e4, 64'h608002f70},{64'h500801018000100, 64'h0, 64'hbf938e117c52b600, 64'h345d19a3ef9367, 64'hbb40051d0011a4, 64'h1a8000000},{64'h6000800000000002, 64'h4014, 64'h43f3462f5c000000, 64'h366000d984a43f, 64'h1e00000549000000, 64'h93ee84b59},{64'h20000041940, 64'h149000000002000, 64'h5ec9ae0000000000, 64'h16400116f4ad6b, 64'h751366000, 64'h199c000000},{64'h418025000000000, 64'h6100, 64'h17960000000000, 64'h31028001a1819000, 64'h99e84d314d3b34, 64'hac57d8000},{64'h2200000000030100, 64'h14, 64'h1f148e2b2c000000, 64'h306ff001d5c63249, 64'h8f1168c0000011e2, 64'h255e},{64'h430003000051000, 64'h1000, 64'hdae217c46f800, 64'hc8ed9816, 64'h6c66ba1b001144, 64'h1767a50000},{64'h1000000000, 64'h200c, 64'h9b60000000000, 64'h12000001cea3501c, 64'h2dd42fa517000ed4, 64'h177c185d56},{64'h5080000000, 64'h4400000000000010, 64'h2794b62abc31a34c, 64'h498000008d80074f, 64'h6380000000107f, 64'hbc0002b10},{64'h400008000100, 64'h0, 64'h29d466117c000000, 64'h4650004f800645, 64'h711000000, 64'h178c000000},{64'h4000010000500c0, 64'h2000, 64'h17a60000000000, 64'h1804006fb, 64'h16fc00253001c44, 64'he24000000},{64'h1100000000, 64'h4280, 64'h0, 64'hd80000119c00000, 64'h150d, 64'h19dcdb8000},{64'h4508006000000000, 64'h4180, 64'h0, 64'ha100000000000000, 64'hceb851ed42a7944e, 64'hc7f7ea49c},{64'h1000000011000, 64'h0, 64'he7c4000000000, 64'h176dd8800, 64'h22b00021c, 64'h0},{64'h400000000010080, 64'hc, 64'h0, 64'heec00749, 64'h7eee8800000000, 64'h70b0},{64'h200000000040040, 64'h180, 64'h0, 64'hf5400037, 64'hc7400000000000, 64'hc14aa8000},{64'h800000000002, 64'h0, 64'hd160000000000000, 64'h461, 64'h2cc7000059000000, 64'h31c6},{64'h10100, 64'h0, 64'ha5b0000000000, 64'h11f0010fc0028d, 64'h0, 64'hc80003160},{64'h4000000140, 64'h6000, 64'h8500000000000, 64'h1d7, 64'h188c, 64'h9b4000000},{64'h1006080000000, 64'h14, 64'h0, 64'haebb600000000000, 64'h23700141f, 64'h14948b1fb0},{64'h10000, 64'h4280, 64'h12488000000000, 64'h3ac00000, 64'hbcc00000000000, 64'h163f418000},{64'h10080, 64'h0, 64'h0, 64'h60c00031, 64'h0, 64'hec6ff5f40},{64'h42800, 64'h0, 64'h9504000000000, 64'ha36b5800, 64'h0, 64'h1a3c000000},{64'h0, 64'h0, 64'h0, 64'h0, 64'h5d1000000, 64'h0},{64'h0, 64'h4000, 64'h0, 64'h0, 64'hbe400000000000, 64'h152c000000},{64'h40, 64'h0, 64'h0, 64'h33, 64'h0, 64'h1a24000000},{64'h4020000, 64'h0, 64'h0, 64'h47900118400000, 64'h1464, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h74b000000, 64'h0},{64'h300000000000002, 64'h4008, 64'h8d60000000000000, 64'h73b, 64'hc400000000000, 64'h12d4007530},{64'h2000000000000000, 64'h10, 64'h0, 64'h237, 64'he200000000000000, 64'h5fd5},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h544000000},{64'h0, 64'h10, 64'h0, 64'h0, 64'h0, 64'h31f0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h150c, 64'h0},{64'h40000, 64'h0, 64'h0, 64'hd9c00000, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'hc7400000000000, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h3210},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'hedc00000, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h5ff0},{64'h0, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0},{64'h1, 64'h0, 64'h0, 64'h0, 64'h0, 64'h0}};

//For 1st BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_A_addr;
reg [63:0]bram_ZYNQ_block_A_din;
wire [63:0]bram_ZYNQ_block_A_dout;
wire bram_ZYNQ_block_A_en;
wire [3:0]bram_ZYNQ_block_A_we;

//For 2nd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_B_addr;
reg [63:0]bram_ZYNQ_block_B_din;
wire [63:0]bram_ZYNQ_block_B_dout;
wire bram_ZYNQ_block_B_en;
wire [3:0]bram_ZYNQ_block_B_we;

//For 3rd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_C_addr;
reg [63:0]bram_ZYNQ_block_C_din;
wire [63:0]bram_ZYNQ_block_C_dout;
wire bram_ZYNQ_block_C_en;
wire [3:0]bram_ZYNQ_block_C_we;

//For 4th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_D_addr;
reg [63:0]bram_ZYNQ_block_D_din;
wire [63:0]bram_ZYNQ_block_D_dout;
wire bram_ZYNQ_block_D_en;
wire [3:0]bram_ZYNQ_block_D_we;

//For 5th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_E_addr;
reg [63:0]bram_ZYNQ_block_E_din;
wire [63:0]bram_ZYNQ_block_E_dout;
wire bram_ZYNQ_block_E_en;
wire [3:0]bram_ZYNQ_block_E_we;

//For 6th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_F_addr;
reg [63:0]bram_ZYNQ_block_F_din;
wire [63:0]bram_ZYNQ_block_F_dout;
wire bram_ZYNQ_block_F_en;
wire [3:0]bram_ZYNQ_block_F_we;

//For 7th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_G_addr;
reg [63:0]bram_ZYNQ_block_G_din;
wire [63:0]bram_ZYNQ_block_G_dout;
wire bram_ZYNQ_block_G_en;
wire [3:0]bram_ZYNQ_block_G_we;

//For 8th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_H_addr;
reg [63:0]bram_ZYNQ_block_H_din;
wire [63:0]bram_ZYNQ_block_H_dout;
wire bram_ZYNQ_block_H_en;
wire [3:0]bram_ZYNQ_block_H_we;

//Instruction BRAM
wire [63:0]bram_ZYNQ_INST_addr;
wire bram_ZYNQ_INST_en;
wire bram_ZYNQ_INST_we;

wire [63:0]bram_ZYNQ_INST_din_part_0;
wire [63:0]bram_ZYNQ_INST_din_part_1;
wire [63:0]bram_ZYNQ_INST_din_part_2;
wire [63:0]bram_ZYNQ_INST_din_part_3;
wire [63:0]bram_ZYNQ_INST_din_part_4;
wire [63:0]bram_ZYNQ_INST_din_part_5;

wire [63:0]bram_ZYNQ_INST_dout_part_0;
wire [63:0]bram_ZYNQ_INST_dout_part_1;
wire [63:0]bram_ZYNQ_INST_dout_part_2;
wire [63:0]bram_ZYNQ_INST_dout_part_3;
wire [63:0]bram_ZYNQ_INST_dout_part_4;
wire [63:0]bram_ZYNQ_INST_dout_part_5;

//debug signals
wire [1:0]debug_state;

reg [31:0]fptr,fptr2;
integer count;
reg complete_bit;

//Mux signals for Address
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_dout;
reg [1:0]sel_mux_dataBRAM;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_dout;

//Mux signals for enable
reg mux_dataBRAM_A_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_en1 = 0; //For clearing
reg mux_dataBRAM_A_en2 = 0; //For loading A matrix
reg mux_dataBRAM_A_en3 = 0; //Currently unused
wire mux_dataBRAM_A_endout;

reg mux_dataBRAM_B_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_en1 = 0; //For clearing
reg mux_dataBRAM_B_en2 = 0; //For loading A matrix
reg mux_dataBRAM_B_en3 = 0; //Currently unused
wire mux_dataBRAM_B_endout;

reg mux_dataBRAM_C_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_en1 = 0; //For clearing
reg mux_dataBRAM_C_en2 = 0; //For loading A matrix
reg mux_dataBRAM_C_en3 = 0; //Currently unused
wire mux_dataBRAM_C_endout;

reg mux_dataBRAM_D_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_en1 = 0; //For clearing
reg mux_dataBRAM_D_en2 = 0; //For loading A matrix
reg mux_dataBRAM_D_en3 = 0; //Currently unused
wire mux_dataBRAM_D_endout;

reg mux_dataBRAM_E_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_E_en1 = 0; //For clearing
reg mux_dataBRAM_E_en2 = 0; //For loading A matrix
reg mux_dataBRAM_E_en3 = 0; //Currently unused
wire mux_dataBRAM_E_endout;

reg mux_dataBRAM_F_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_F_en1 = 0; //For clearing
reg mux_dataBRAM_F_en2 = 0; //For loading A matrix
reg mux_dataBRAM_F_en3 = 0; //Currently unused
wire mux_dataBRAM_F_endout;

reg mux_dataBRAM_G_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_G_en1 = 0; //For clearing
reg mux_dataBRAM_G_en2 = 0; //For loading A matrix
reg mux_dataBRAM_G_en3 = 0; //Currently unused
wire mux_dataBRAM_G_endout;

reg mux_dataBRAM_H_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_H_en1 = 0; //For clearing
reg mux_dataBRAM_H_en2 = 0; //For loading A matrix
reg mux_dataBRAM_H_en3 = 0; //Currently unused
wire mux_dataBRAM_H_endout;

//Mux signals for write enable
reg mux_dataBRAM_A_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_we1 = 0; //For clearing
reg mux_dataBRAM_A_we2 = 0; //For loading A matrix
reg mux_dataBRAM_A_we3 = 0; //Currently unused
wire mux_dataBRAM_A_wedout;

reg mux_dataBRAM_B_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_we1 = 0; //For clearing
reg mux_dataBRAM_B_we2 = 0; //For loading A matrix
reg mux_dataBRAM_B_we3 = 0; //Currently unused
wire mux_dataBRAM_B_wedout;

reg mux_dataBRAM_C_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_we1 = 0; //For clearing
reg mux_dataBRAM_C_we2 = 0; //For loading A matrix
reg mux_dataBRAM_C_we3 = 0; //Currently unused
wire mux_dataBRAM_C_wedout;

reg mux_dataBRAM_D_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_we1 = 0; //For clearing
reg mux_dataBRAM_D_we2 = 0; //For loading A matrix
reg mux_dataBRAM_D_we3 = 0; //Currently unused
wire mux_dataBRAM_D_wedout;

reg mux_dataBRAM_E_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_E_we1 = 0; //For clearing
reg mux_dataBRAM_E_we2 = 0; //For loading A matrix
reg mux_dataBRAM_E_we3 = 0; //Currently unused
wire mux_dataBRAM_E_wedout;

reg mux_dataBRAM_F_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_F_we1 = 0; //For clearing
reg mux_dataBRAM_F_we2 = 0; //For loading A matrix
reg mux_dataBRAM_F_we3 = 0; //Currently unused
wire mux_dataBRAM_F_wedout;

reg mux_dataBRAM_G_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_G_we1 = 0; //For clearing
reg mux_dataBRAM_G_we2 = 0; //For loading A matrix
reg mux_dataBRAM_G_we3 = 0; //Currently unused
wire mux_dataBRAM_G_wedout;

reg mux_dataBRAM_H_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_H_we1 = 0; //For clearing
reg mux_dataBRAM_H_we2 = 0; //For loading A matrix
reg mux_dataBRAM_H_we3 = 0; //Currently unused
wire mux_dataBRAM_H_wedout;

//Mux signals for din
reg [63:0]mux_dataBRAM_A_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_A_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_A_din_out;
reg sel_mux_dataBRAM_din;

reg [63:0]mux_dataBRAM_B_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_B_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_B_din_out;

reg [63:0]mux_dataBRAM_C_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_C_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_C_din_out;

reg [63:0]mux_dataBRAM_D_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_D_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_D_din_out;

reg [63:0]mux_dataBRAM_E_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_E_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_E_din_out;

reg [63:0]mux_dataBRAM_F_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_F_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_F_din_out;

reg [63:0]mux_dataBRAM_G_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_G_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_G_din_out;

reg [63:0]mux_dataBRAM_H_din0; //for clearing the data BRAMS
reg [63:0]mux_dataBRAM_H_din1; //for loading the data BRAMS
wire [63:0]mux_dataBRAM_H_din_out;

//Instruction BRAM muxes
reg [63:0]instBRAM_part0_din;
reg [63:0]instBRAM_part1_din;
reg [63:0]instBRAM_part2_din;
reg [63:0]instBRAM_part3_din;
reg [63:0]instBRAM_part4_din;
reg [63:0]instBRAM_part5_din;

reg instBRAM_en = 0;
reg instBRAM_we = 0;
reg [ADDR_WIDTH-1:0]instBRAM_addr;


//Memory dump start and complete signals
reg start_mem_dump;
reg mem_dump_complete;
reg start_dataBRAM_erase;
reg dataBRAM_erase_complete;
reg start_A_load;
reg A_load_complete;
reg start_instBRAM_erase;
reg instBRAM_erase_complete;
reg start_inst_load;
reg inst_load_complete;
reg start_full_run;
reg complete_full_run;
reg start0; //For full run
reg complete_sig;

LUDH_TEST_WRAPPER #(ADDR_WIDTH,ADDR_WIDTH_DATA_BRAM,CTRL_WIDTH,AU_SEL_WIDTH,BRAM_SEL_WIDTH) uut1 (
CLK_100,

locked,
RST_IN,
start_sig,
completed,

//First BRAM
bram_ZYNQ_block_A_addr, 
bram_ZYNQ_block_A_din, 
bram_ZYNQ_block_A_dout, 
bram_ZYNQ_block_A_en,
bram_ZYNQ_block_A_we, 

//Second BRAM
bram_ZYNQ_block_B_addr, 
bram_ZYNQ_block_B_din, 
bram_ZYNQ_block_B_dout, 
bram_ZYNQ_block_B_en,
bram_ZYNQ_block_B_we, 

//Third BRAM
bram_ZYNQ_block_C_addr, 
bram_ZYNQ_block_C_din, 
bram_ZYNQ_block_C_dout, 
bram_ZYNQ_block_C_en,
bram_ZYNQ_block_C_we, 

//Fourth BRAM
bram_ZYNQ_block_D_addr, 
bram_ZYNQ_block_D_din, 
bram_ZYNQ_block_D_dout, 
bram_ZYNQ_block_D_en,
bram_ZYNQ_block_D_we, 

//Fifth BRAM
bram_ZYNQ_block_E_addr, 
bram_ZYNQ_block_E_din, 
bram_ZYNQ_block_E_dout, 
bram_ZYNQ_block_E_en,
bram_ZYNQ_block_E_we, 

//Sixth BRAM
bram_ZYNQ_block_F_addr, 
bram_ZYNQ_block_F_din, 
bram_ZYNQ_block_F_dout, 
bram_ZYNQ_block_F_en,
bram_ZYNQ_block_F_we, 

//Seventh BRAM
bram_ZYNQ_block_G_addr, 
bram_ZYNQ_block_G_din, 
bram_ZYNQ_block_G_dout, 
bram_ZYNQ_block_G_en,
bram_ZYNQ_block_G_we, 

//Eighth BRAM
bram_ZYNQ_block_H_addr, 
bram_ZYNQ_block_H_din, 
bram_ZYNQ_block_H_dout, 
bram_ZYNQ_block_H_en,
bram_ZYNQ_block_H_we, 

//Instruction BRAM
bram_ZYNQ_INST_addr,
bram_ZYNQ_INST_en,
bram_ZYNQ_INST_we,
        
bram_ZYNQ_INST_din_part_0,
bram_ZYNQ_INST_din_part_1,
bram_ZYNQ_INST_din_part_2,
bram_ZYNQ_INST_din_part_3,
bram_ZYNQ_INST_din_part_4,
bram_ZYNQ_INST_din_part_5,
        
bram_ZYNQ_INST_dout_part_0,
bram_ZYNQ_INST_dout_part_1,
bram_ZYNQ_INST_dout_part_2,
bram_ZYNQ_INST_dout_part_3,
bram_ZYNQ_INST_dout_part_4,
bram_ZYNQ_INST_dout_part_5,
        
//debug signals
debug_state
);

initial begin
CLK_100 = 1'b1;
forever #(t_100/2) CLK_100 = ~CLK_100;
end

//Initiallizing the mux to be used for DATA BRAMS address multiplexing
//For address
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut2(mux_dataBRAM_A_dout,mux_dataBRAM_A_0,mux_dataBRAM_A_1,mux_dataBRAM_A_2,mux_dataBRAM_A_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut3(mux_dataBRAM_B_dout,mux_dataBRAM_B_0,mux_dataBRAM_B_1,mux_dataBRAM_B_2,mux_dataBRAM_B_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut4(mux_dataBRAM_C_dout,mux_dataBRAM_C_0,mux_dataBRAM_C_1,mux_dataBRAM_C_2,mux_dataBRAM_C_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut5(mux_dataBRAM_D_dout,mux_dataBRAM_D_0,mux_dataBRAM_D_1,mux_dataBRAM_D_2,mux_dataBRAM_D_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut18(mux_dataBRAM_E_dout,mux_dataBRAM_E_0,mux_dataBRAM_E_1,mux_dataBRAM_E_2,mux_dataBRAM_E_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut19(mux_dataBRAM_F_dout,mux_dataBRAM_F_0,mux_dataBRAM_F_1,mux_dataBRAM_F_2,mux_dataBRAM_F_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut20(mux_dataBRAM_G_dout,mux_dataBRAM_G_0,mux_dataBRAM_G_1,mux_dataBRAM_G_2,mux_dataBRAM_G_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut21(mux_dataBRAM_H_dout,mux_dataBRAM_H_0,mux_dataBRAM_H_1,mux_dataBRAM_H_2,mux_dataBRAM_H_3,sel_mux_dataBRAM);

//For enable
mux_4x1 #(1) uut6(mux_dataBRAM_A_endout,mux_dataBRAM_A_en0,mux_dataBRAM_A_en1,mux_dataBRAM_A_en2,mux_dataBRAM_A_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut7(mux_dataBRAM_B_endout,mux_dataBRAM_B_en0,mux_dataBRAM_B_en1,mux_dataBRAM_B_en2,mux_dataBRAM_B_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut8(mux_dataBRAM_C_endout,mux_dataBRAM_C_en0,mux_dataBRAM_C_en1,mux_dataBRAM_C_en2,mux_dataBRAM_C_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut9(mux_dataBRAM_D_endout,mux_dataBRAM_D_en0,mux_dataBRAM_D_en1,mux_dataBRAM_D_en2,mux_dataBRAM_D_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut22(mux_dataBRAM_E_endout,mux_dataBRAM_E_en0,mux_dataBRAM_E_en1,mux_dataBRAM_E_en2,mux_dataBRAM_E_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut23(mux_dataBRAM_F_endout,mux_dataBRAM_F_en0,mux_dataBRAM_F_en1,mux_dataBRAM_F_en2,mux_dataBRAM_F_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut24(mux_dataBRAM_G_endout,mux_dataBRAM_G_en0,mux_dataBRAM_G_en1,mux_dataBRAM_G_en2,mux_dataBRAM_G_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut25(mux_dataBRAM_H_endout,mux_dataBRAM_H_en0,mux_dataBRAM_H_en1,mux_dataBRAM_H_en2,mux_dataBRAM_H_en3,sel_mux_dataBRAM);

//For Write enable
mux_4x1 #(1) uut10(mux_dataBRAM_A_wedout,mux_dataBRAM_A_we0,mux_dataBRAM_A_we1,mux_dataBRAM_A_we2,mux_dataBRAM_A_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut11(mux_dataBRAM_B_wedout,mux_dataBRAM_B_we0,mux_dataBRAM_B_we1,mux_dataBRAM_B_we2,mux_dataBRAM_B_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut12(mux_dataBRAM_C_wedout,mux_dataBRAM_C_we0,mux_dataBRAM_C_we1,mux_dataBRAM_C_we2,mux_dataBRAM_C_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut13(mux_dataBRAM_D_wedout,mux_dataBRAM_D_we0,mux_dataBRAM_D_we1,mux_dataBRAM_D_we2,mux_dataBRAM_D_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut26(mux_dataBRAM_E_wedout,mux_dataBRAM_E_we0,mux_dataBRAM_E_we1,mux_dataBRAM_E_we2,mux_dataBRAM_E_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut27(mux_dataBRAM_F_wedout,mux_dataBRAM_F_we0,mux_dataBRAM_F_we1,mux_dataBRAM_F_we2,mux_dataBRAM_F_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut28(mux_dataBRAM_G_wedout,mux_dataBRAM_G_we0,mux_dataBRAM_G_we1,mux_dataBRAM_G_we2,mux_dataBRAM_G_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut29(mux_dataBRAM_H_wedout,mux_dataBRAM_H_we0,mux_dataBRAM_H_we1,mux_dataBRAM_H_we2,mux_dataBRAM_H_we3,sel_mux_dataBRAM);

//For din
mux_2x1 #(64) uut14(mux_dataBRAM_A_din_out,mux_dataBRAM_A_din0,mux_dataBRAM_A_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut15(mux_dataBRAM_B_din_out,mux_dataBRAM_B_din0,mux_dataBRAM_B_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut16(mux_dataBRAM_C_din_out,mux_dataBRAM_C_din0,mux_dataBRAM_C_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut17(mux_dataBRAM_D_din_out,mux_dataBRAM_D_din0,mux_dataBRAM_D_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut30(mux_dataBRAM_E_din_out,mux_dataBRAM_E_din0,mux_dataBRAM_E_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut31(mux_dataBRAM_F_din_out,mux_dataBRAM_F_din0,mux_dataBRAM_F_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut32(mux_dataBRAM_G_din_out,mux_dataBRAM_G_din0,mux_dataBRAM_G_din1,sel_mux_dataBRAM_din);
mux_2x1 #(64) uut33(mux_dataBRAM_H_din_out,mux_dataBRAM_H_din0,mux_dataBRAM_H_din1,sel_mux_dataBRAM_din);


initial begin
start_mem_dump <= 0;
mem_dump_complete <= 0;
start_dataBRAM_erase <= 0;
dataBRAM_erase_complete <= 0;
start_A_load <= 0;
A_load_complete <= 0;
start_instBRAM_erase <= 0;
instBRAM_erase_complete <= 0;
start_inst_load <= 0;
inst_load_complete <= 0;
complete_full_run <= 0;
sel_mux_dataBRAM <= 2'b00;
sel_mux_dataBRAM_din <= 1'b0;

count <= -1;
complete_bit <= 1'b0;
locked <= 1'b0;

#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
RST_IN <= 1'b1;

//Resetting the contents of data BRAMS and Inst BRAM
#(t_100*50)
sel_mux_dataBRAM <= 2'b01;
sel_mux_dataBRAM_din <= 1'b0;
start_dataBRAM_erase <= 1'b1;

@(posedge dataBRAM_erase_complete)
#(t_100*50)
start_dataBRAM_erase <= 0;

#(t_100*50)
start_instBRAM_erase <= 1'b1;

@(posedge instBRAM_erase_complete)
#(t_100*50)
start_instBRAM_erase <= 0;

//Loading the A matrix
#(t_100*50)
sel_mux_dataBRAM <= 2'b10;
sel_mux_dataBRAM_din <= 1'b1;
start_A_load <= 1'b1;

@(posedge A_load_complete)
#(t_100*50)
start_A_load <= 0;

//RST = 0
#(t_100*50)
RST_IN <= 1'b0;

//Locked = 1
#(t_100*50)
locked <= 1'b1;

//Loading the instruction matrix and starting LU Decomposition
#(t_100*50)
start_full_run = 1'b1;

@(posedge complete_sig)
complete_bit <= 1'b1;
#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
sel_mux_dataBRAM <= 2'b00;
start_mem_dump <= 1;

@(posedge mem_dump_complete)
#(t_100*50)
start_mem_dump <= 0;
$stop;

end

assign start_sig = start0;
assign complete_sig = complete_full_run;

//Address signals(data BRAM)
assign bram_ZYNQ_block_A_addr = mux_dataBRAM_A_dout;
assign bram_ZYNQ_block_B_addr = mux_dataBRAM_B_dout;
assign bram_ZYNQ_block_C_addr = mux_dataBRAM_C_dout;
assign bram_ZYNQ_block_D_addr = mux_dataBRAM_D_dout;
assign bram_ZYNQ_block_E_addr = mux_dataBRAM_E_dout;
assign bram_ZYNQ_block_F_addr = mux_dataBRAM_F_dout;
assign bram_ZYNQ_block_G_addr = mux_dataBRAM_G_dout;
assign bram_ZYNQ_block_H_addr = mux_dataBRAM_H_dout;

//Enable signals(data BRAM)
assign bram_ZYNQ_block_A_en = mux_dataBRAM_A_endout;
assign bram_ZYNQ_block_B_en = mux_dataBRAM_B_endout;
assign bram_ZYNQ_block_C_en = mux_dataBRAM_C_endout;
assign bram_ZYNQ_block_D_en = mux_dataBRAM_D_endout;
assign bram_ZYNQ_block_E_en = mux_dataBRAM_E_endout;
assign bram_ZYNQ_block_F_en = mux_dataBRAM_F_endout;
assign bram_ZYNQ_block_G_en = mux_dataBRAM_G_endout;
assign bram_ZYNQ_block_H_en = mux_dataBRAM_H_endout;

//Write enable signals(data BRAM)
assign bram_ZYNQ_block_A_we = mux_dataBRAM_A_wedout;
assign bram_ZYNQ_block_B_we = mux_dataBRAM_B_wedout;
assign bram_ZYNQ_block_C_we = mux_dataBRAM_C_wedout;
assign bram_ZYNQ_block_D_we = mux_dataBRAM_D_wedout;
assign bram_ZYNQ_block_E_we = mux_dataBRAM_E_wedout;
assign bram_ZYNQ_block_F_we = mux_dataBRAM_F_wedout;
assign bram_ZYNQ_block_G_we = mux_dataBRAM_G_wedout;
assign bram_ZYNQ_block_H_we = mux_dataBRAM_H_wedout;

//din signals(data BRAM)
assign bram_ZYNQ_block_A_din = mux_dataBRAM_A_din_out;
assign bram_ZYNQ_block_B_din = mux_dataBRAM_B_din_out;
assign bram_ZYNQ_block_C_din = mux_dataBRAM_C_din_out;
assign bram_ZYNQ_block_D_din = mux_dataBRAM_D_din_out;
assign bram_ZYNQ_block_E_din = mux_dataBRAM_E_din_out;
assign bram_ZYNQ_block_F_din = mux_dataBRAM_F_din_out;
assign bram_ZYNQ_block_G_din = mux_dataBRAM_G_din_out;
assign bram_ZYNQ_block_H_din = mux_dataBRAM_H_din_out;

//Address signal(inst BRAM)
assign bram_ZYNQ_INST_addr = instBRAM_addr;

//Enable signal(inst BRAM)
assign bram_ZYNQ_INST_en = instBRAM_en;

//Write enable signal(inst BRAM)
assign bram_ZYNQ_INST_we = instBRAM_we;

//din signal(inst BRAM)
assign bram_ZYNQ_INST_din_part_0 = instBRAM_part0_din;
assign bram_ZYNQ_INST_din_part_1 = instBRAM_part1_din;
assign bram_ZYNQ_INST_din_part_2 = instBRAM_part2_din;
assign bram_ZYNQ_INST_din_part_3 = instBRAM_part3_din;
assign bram_ZYNQ_INST_din_part_4 = instBRAM_part4_din;
assign bram_ZYNQ_INST_din_part_5 = instBRAM_part5_din;


//Always block for full run
always@(posedge CLK_100) begin
if(CLK_100  == 1 && start_full_run == 1 && complete_full_run != 1) begin
//Start loading complete instructions
start_inst_load <= 1'b1;
@(posedge inst_load_complete)
#(t_100*50)
start_inst_load <= 0;

//Start the LU Decomposition
#(t_100*50)
start0 <= 1'b1;
complete_full_run <= 1'b0;

//Waiting for completion
@(posedge completed)
complete_full_run <= 1'b1;

end
else if(CLK_100 == 1 && start_full_run == 0) begin
start0 <= 0;
complete_full_run <= 0;
end
end

//Always block to dump bram contents
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_mem_dump == 1 && mem_dump_complete != 1)begin 

    if(count == -1) begin
        fptr = $fopen("BRAM_dump.txt","w");
        $fdisplay(fptr,"float bram_dump[%d][%d];",BRAM_LIMIT_IND_DEBUG,DATA_BRAM_SIZE);
        mux_dataBRAM_A_en0 = 1'b1; mux_dataBRAM_B_en0 = 1'b1; mux_dataBRAM_C_en0 = 1'b1; mux_dataBRAM_D_en0 = 1'b1; mux_dataBRAM_E_en0 = 1'b1; mux_dataBRAM_F_en0 = 1'b1; mux_dataBRAM_G_en0 = 1'b1; mux_dataBRAM_H_en0 = 1'b1;
        mux_dataBRAM_A_we0 = 1'b0; mux_dataBRAM_B_we0 = 1'b0; mux_dataBRAM_C_we0 = 1'b0; mux_dataBRAM_D_we0 = 1'b0; mux_dataBRAM_E_we0 = 1'b0; mux_dataBRAM_F_we0 = 1'b0; mux_dataBRAM_G_we0 = 1'b0; mux_dataBRAM_H_we0 = 1'b0;
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];
    end
    else if(count == 0) begin
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Addres
    end
    else if(count <= DATA_BRAM_SIZE && count >= 1)begin
        $fdisplay(fptr,"bram_dump[0][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_A_dout)); //count-1 because BRAM has single cycle latency
        $fdisplay(fptr,"bram_dump[1][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_B_dout));
        $fdisplay(fptr,"bram_dump[2][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_C_dout));
        $fdisplay(fptr,"bram_dump[3][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_D_dout));
        $fdisplay(fptr,"bram_dump[4][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_E_dout));
        $fdisplay(fptr,"bram_dump[5][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_F_dout));
        $fdisplay(fptr,"bram_dump[6][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_G_dout));
        $fdisplay(fptr,"bram_dump[7][%d] = %1.17e;",count-1,float_conv(bram_ZYNQ_block_H_dout));
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Address
    end
    else if (count == DATA_BRAM_SIZE+1) begin
        $fclose(fptr);
        count = -1;
        mem_dump_complete = 1;    
        mux_dataBRAM_A_en0 = 1'b0; mux_dataBRAM_B_en0 = 1'b0; mux_dataBRAM_C_en0 = 1'b0; mux_dataBRAM_D_en0 = 1'b0; mux_dataBRAM_E_en0 = 1'b0; mux_dataBRAM_F_en0 = 1'b0; mux_dataBRAM_G_en0 = 1'b0; mux_dataBRAM_H_en0 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_mem_dump == 0)
    mem_dump_complete = 0;
end


//Always block to erase data BRAM contents
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_dataBRAM_erase == 1 && dataBRAM_erase_complete != 1)begin 

    if(count <= DATA_BRAM_SIZE-2 && count >= -1)begin
        if(count == -1) begin
            mux_dataBRAM_A_en1 = 1'b1; mux_dataBRAM_B_en1 = 1'b1; mux_dataBRAM_C_en1 = 1'b1; mux_dataBRAM_D_en1 = 1'b1; mux_dataBRAM_E_en1 = 1'b1; mux_dataBRAM_F_en1 = 1'b1; mux_dataBRAM_G_en1 = 1'b1; mux_dataBRAM_H_en1 = 1'b1;
            mux_dataBRAM_A_we1 = 1'b1; mux_dataBRAM_B_we1 = 1'b1; mux_dataBRAM_C_we1 = 1'b1; mux_dataBRAM_D_we1 = 1'b1; mux_dataBRAM_E_we1 = 1'b1; mux_dataBRAM_F_we1 = 1'b1; mux_dataBRAM_G_we1 = 1'b1; mux_dataBRAM_H_we1 = 1'b1;
            mux_dataBRAM_A_din0 = 0; mux_dataBRAM_B_din0 = 0; mux_dataBRAM_C_din0 = 0; mux_dataBRAM_D_din0 = 0; mux_dataBRAM_E_din0 = 0; mux_dataBRAM_F_din0 = 0; mux_dataBRAM_G_din0 = 0; mux_dataBRAM_H_din0 = 0; //Reset value
        end
        count = count + 1;
        mux_dataBRAM_A_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; //Address
    end
    else if (count == DATA_BRAM_SIZE-1) begin
        count = -1;
        dataBRAM_erase_complete = 1;   
        mux_dataBRAM_A_en1 = 1'b0; mux_dataBRAM_B_en1 = 1'b0; mux_dataBRAM_C_en1 = 1'b0; mux_dataBRAM_D_en1 = 1'b0; mux_dataBRAM_E_en1 = 1'b0; mux_dataBRAM_F_en1 = 1'b0; mux_dataBRAM_G_en1 = 1'b0; mux_dataBRAM_H_en1 = 1'b0;
        mux_dataBRAM_A_we1 = 1'b0; mux_dataBRAM_B_we1 = 1'b0; mux_dataBRAM_C_we1 = 1'b0; mux_dataBRAM_D_we1 = 1'b0; mux_dataBRAM_E_we1 = 1'b0; mux_dataBRAM_F_we1 = 1'b0; mux_dataBRAM_G_we1 = 1'b0; mux_dataBRAM_H_we1 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_dataBRAM_erase == 0)
    dataBRAM_erase_complete = 0;
end

//Always block to load the A matrix in data bram
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_A_load == 1 && A_load_complete != 1)begin 

    if(count <= A_size-2 && count >= -1)begin
        if(count == -1) //Initialization of en signals
            mux_dataBRAM_A_en2 = 1'b1; mux_dataBRAM_B_en2 = 1'b1; mux_dataBRAM_C_en2 = 1'b1; mux_dataBRAM_D_en2 = 1'b1; mux_dataBRAM_E_en2 = 1'b1; mux_dataBRAM_F_en2 = 1'b1; mux_dataBRAM_G_en2 = 1'b1; mux_dataBRAM_H_en2 = 1'b1;
            
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0; mux_dataBRAM_E_we2 = 1'b0; mux_dataBRAM_F_we2 = 1'b0; mux_dataBRAM_G_we2 = 1'b0; mux_dataBRAM_H_we2 = 1'b0;//Initially assigning all the write enables to 0
        count = count + 1;
        if(A_BRAMInd[count] == 0) begin//making one of the write enables 1
            mux_dataBRAM_A_we2 = 1'b1; mux_dataBRAM_A_2 = A_BRAMAddr[count]; mux_dataBRAM_A_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 1) begin
            mux_dataBRAM_B_we2 = 1'b1; mux_dataBRAM_B_2 = A_BRAMAddr[count]; mux_dataBRAM_B_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 2) begin
            mux_dataBRAM_C_we2 = 1'b1; mux_dataBRAM_C_2 = A_BRAMAddr[count]; mux_dataBRAM_C_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 3) begin
            mux_dataBRAM_D_we2 = 1'b1; mux_dataBRAM_D_2 = A_BRAMAddr[count]; mux_dataBRAM_D_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 4) begin
            mux_dataBRAM_E_we2 = 1'b1; mux_dataBRAM_E_2 = A_BRAMAddr[count]; mux_dataBRAM_E_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 5) begin
            mux_dataBRAM_F_we2 = 1'b1; mux_dataBRAM_F_2 = A_BRAMAddr[count]; mux_dataBRAM_F_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 6) begin
            mux_dataBRAM_G_we2 = 1'b1; mux_dataBRAM_G_2 = A_BRAMAddr[count]; mux_dataBRAM_G_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 7) begin
            mux_dataBRAM_H_we2 = 1'b1; mux_dataBRAM_H_2 = A_BRAMAddr[count]; mux_dataBRAM_H_din1 = A[count];
        end
    end
    else if (count == A_size-1) begin
        count = -1;
        A_load_complete = 1;   
        mux_dataBRAM_A_en2 = 1'b0; mux_dataBRAM_B_en2 = 1'b0; mux_dataBRAM_C_en2 = 1'b0; mux_dataBRAM_D_en2 = 1'b0; mux_dataBRAM_E_en2 = 1'b0; mux_dataBRAM_F_en2 = 1'b0; mux_dataBRAM_G_en2 = 1'b0; mux_dataBRAM_H_en2 = 1'b0;
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0; mux_dataBRAM_E_we2 = 1'b0; mux_dataBRAM_F_we2 = 1'b0; mux_dataBRAM_G_we2 = 1'b0; mux_dataBRAM_H_we2 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_A_load == 0)
    A_load_complete = 0;
end

//Always block to erase inst BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_instBRAM_erase == 1 && instBRAM_erase_complete != 1)begin 

    if(count <= INST_BRAM_SIZE-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
            instBRAM_part0_din = 0; instBRAM_part1_din = 0; instBRAM_part2_din = 0; instBRAM_part3_din = 0; instBRAM_part4_din = 0; instBRAM_part5_din = 0;
        end
        count = count + 1;
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == INST_BRAM_SIZE-1) begin
        count = -1;
        instBRAM_erase_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_instBRAM_erase == 0)
    instBRAM_erase_complete = 0;
end

//Always block to load instruction to instruction BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_inst_load == 1 && inst_load_complete != 1)begin 

    if(count <= total_instructions-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
        end
        count = count + 1;
        instBRAM_part0_din = Inst[count][0]; instBRAM_part1_din = Inst[count][1]; instBRAM_part2_din = Inst[count][2]; instBRAM_part3_din = Inst[count][3]; 
        instBRAM_part4_din = Inst[count][4]; instBRAM_part5_din = Inst[count][5];
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == total_instructions-1) begin
        count = -1;
        inst_load_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_inst_load == 0)
    inst_load_complete = 0;
end

function real float_conv(input [63:0]b_num);
reg sign;
reg [10:0]weighted_expt;
integer actual_expt;
reg [1:52] mantissa;
reg [10:0] i;
static real real_one = 1.0;
static longint long_one = 1;
real temp_result,temp_decimal;

begin
sign = b_num >> 63;
weighted_expt = (b_num & 64'h7ff0000000000000)>> 52;
mantissa = b_num & 64'h000fffffffffffff;
if(weighted_expt == 0)begin
	temp_result = 1.0;
	for(i=0;i<1022;i=i+1)
		temp_result = temp_result/2;

	temp_decimal = 0;
	for(i=1;i<=52;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(real_one/(long_one<<i));
		
	temp_result = temp_result*temp_decimal;
	if(sign==1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
	end
else if(weighted_expt>0 && weighted_expt <2047) begin
	actual_expt = weighted_expt-1023;
	if(actual_expt<0)begin
		temp_result = 1.0;
		actual_expt = -actual_expt;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result/2;
		end
	else begin
		temp_result = 1.0;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result*2;
	end

	temp_decimal = 0;
	for(i=1;i<=52;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(real_one/(long_one<<i));

	temp_decimal = temp_decimal + 1;
	temp_result = temp_result*temp_decimal;
	if(sign == 1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
end
else if(weighted_expt == 2047)begin
/*if(mantissa == 0 and sign == 0)
float_conv = "inf";
else if(mantissa == 0 and sign == 1)
float_conv = "-inf";
else
float_conv = "nan";*/
end

end
endfunction

endmodule

module mux_4x1 #(parameter integer data_width = 11)(dout,din0,din1,din2,din3,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input [data_width-1:0]din2;
input [data_width-1:0]din3;
input [1:0]sel;

always@(din0,din1,din2,din3,sel) begin
case(sel)
2'b00: dout <= din0;
2'b01: dout <= din1;
2'b10: dout <= din2;
2'b11: dout <= din3;
endcase
end
endmodule

module mux_2x1 #(parameter integer data_width = 32)(dout,din0,din1,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input sel;

always@(din0,din1,sel) begin
case(sel)
1'b0: dout <= din0;
1'b1: dout <= din1;
endcase
end
endmodule













