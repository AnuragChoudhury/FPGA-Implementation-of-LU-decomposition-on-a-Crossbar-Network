`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.12.2019 07:59:36
// Design Name: 
// Module Name: simTester_verilog
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simTester_verilog();
reg CLK_100, locked, RST_IN,start_sig;
wire  completed;
localparam time t_100 = 40;

localparam integer ADDR_WIDTH = 12;
localparam integer INST_BRAM_SIZE = 4096;//(2**ADDR_WIDTH)
localparam integer ADDR_WIDTH_DATA_BRAM = 10;
localparam integer DATA_BRAM_SIZE = 1024;//(2**ADDR_WIDTH_DATA_BRAM)
localparam integer CTRL_WIDTH = 357;
localparam integer AU_SEL_WIDTH = 5;
localparam integer BRAM_SEL_WIDTH = 5;

//This parameter = no. of BRAMS
localparam integer BRAM_LIMIT_IND_DEBUG = 8; //It indicates that BRAM contents from location 0 to BRAM_LIMIT_IND_DEBUG will be dumped for all 8 BRAMS for every cycle

//Constant array to load the A matrix
localparam integer A_size = 665;
localparam integer A[0:664] = '{1040747617, -1115125579, -1217732213, -1115125579, 1040747617, -1115125579, -1217732213, -1115125579, 1040747214, -1115125579, -1115125579, -1224329283, 1097859611, -1174758381, -1249495107, -1214841163, -1214841163, -1174724021, 992423598, -1195864924, -1165849545, -1165909675, -1115125579, -1115125579, 906377149, 957052394, 1051382526, -1183765464, -1102263091, -1184933695, -1217732213, -1215940675, -1162860248, 967674385, 1011997911, -1136386606, 961931477, 1040748556, -1115125579, -1208793849, -1115125579, 1040747483, -1115125579, -1115125579, -1218831725, 1089471840, -1172709145, -1249495107, -1206452555, -1207277189, -1172657605, 998327567, -1171437834, -1160343397, -1165325559, -1115125579, -1115125579, 914765757, 961038124, 1051387090, -1177404081, -1102263091, -1183215709, -1208793849, -1205902800, -1150782263, 963030989, 1020614689, -1127997998, 984159544, 1040747617, -1217732213, -1115125579, 1040747214, -1115125579, -1223229771, 1022608091, -1199580608, -1249495107, -1124941055, -1199580608, -1217732213, -1197101875, 1013540878, 944879383, -1215390919, -1156498864, -1115125579, -1115125579, 919163804, -1217732213, 1051372829, 897988541, -1219931236, -1124941055, -1214841163, 1063054788, -1214841163, -1084926640, 1024661085, -1127997998, -1136386606, 1040748556, -1115125579, -1115125579, -1208793849, 1065353216, -1115125579, 1040747483, -1115125579, -1218831725, -1115125579, -1102263091, -1115125579, 1051373332, -1230518868, -1207277189, 916964780, -1208793849, -1127997998, 897988541, 1019532357, -1249495107, -1207002311, -1211542628, -1207552067, -1214291408, 999040532, -1148516131, 932092729, -1207002311, -1148516131, 1054312835, -1209893361, -1093315231, -1127997998, -1218831725, -1241106499, -1209893361, 1019508198, -1223229771, -1202604265, -1156700728, -1198613703, -1213741652, -1136386606, 1013582754, 1065353216, 1040747617, -1217732213, -1115125579, -1217732213, 1011130328, -1215940675, 1040747080, -1115125579, -1228319844, 1003930352, -1223229771, -1222130260, -1143594098, -1115125579, -1115125579, -1214291408, 1051372829, -1228319844, -1222130260, 1011129254, -1217732213, -1136386606, -1084926640, -1215940675, -1143594098, -1217732213, 1062667150, 1074091348, -1084926640, 1065353216, -1093315231, -1084926640, -1115125579, 1040748556, -1115125579, -1208793849, -1115125579, 1040747818, -1115125579, -1214841163, -1102263091, -1115125579, -1115125579, 1051373433, -1210443117, 930850946, -1210443117, -1127997998, -1208793849, 954367503, 1020254449, -1190087656, -1162911788, -1206727433, -1228319844, -1192703828, 1016038938, -1192703828, -1131567116, -1214841163, -1190087656, -1163830911, -1193528462, 1020305988, -1206452555, -1127997998, -1093315231, -1206452555, -1131567116, -1206452555, 1054751022, 1019485650, -1136386606, -1136386606, 1040747617, -1217732213, -1115125579, -1136386606, -1217732213, 1011130328, -1215940675, 1040747080, -1226120821, -1115125579, 1003908877, -1241106499, -1215940675, -1143615573, -1226120821, 1011120664, -1241106499, -1217732213, -1136386606, -1115125579, -1115125579, -1214291408, 1051372829, -1084926640, -1215940675, -1143615573, -1217732213, 1062666999, 1040747617, -1217732213, -1115125579, 1040747214, -1115125579, -1223229771, 1022372941, -1198063947, -1241106499, -1125189627, -1197926508, -1217732213, -1193528462, 1013547320, 945429139, -1216632702, -1156571879, -1115125579, -1115125579, 919163804, -1216632702, 1051372829, 910775196, -1219931236, 1040747617, -1217732213, -1115125579, -1217732213, 1011130328, -1215940675, 1040747080, -1115125579, -1228319844, 1003928204, -1222130260, -1223229771, -1143594098, -1115125579, -1115125579, -1214291408, 1051372829, -1228319844, -1223229771, 1011128180, -1217732213, -1136386606, -1215940675, -1143594098, -1217732213, 1062667150, -1084926640, 1065353216, 1040747617, -1217732213, -1115125579, -1217732213, 1011130328, -1215940675, 1003923909, -1214291408, -1143600541, 1040747080, -1115125579, -1226120821, -1115125579, -1214291408, -1115125579, 1051372829, -1226120821, 1011118516, -1136386606, -1217732213, -1136386606, 1019485650, -1136386606, -1084926640, -1215940675, -1143600541, -1217732213, 1062667100, -1084926640, 1074091348, -1084926640, 1065353216, -1093315231, -1115125579, 1040748556, -1115125579, -1208793849, -1115125579, 1040747818, -1115125579, -1214841163, -1102263091, -1115125579, -1115125579, 1051373433, -1208793849, 930850946, -1212092384, -1127997998, -1208793849, 954230064, 1020251764, -1190087656, -1162963327, -1206727433, -1228319844, -1192841267, 1016011558, -1192703828, -1131594497, -1214841163, -1190087656, -1163899630, -1193665901, 1020301157, -1206452555, -1127997998, -1093315231, -1206452555, -1131594497, -1206452555, 1054749311, -1136386606, -1127997998, 1063159478, -1084926640, 1040747348, -1115125579, -1221030748, 1040747080, -1115125579, -1226120821, -1115125579, -1115125579, 1051372561, -1222130260, -1222130260, 997453004, -1150073593, 897988541, -1249495107, -1150073593, 1062619872, -1215390919, -1215390919, -1084926640, -1226120821, -1215390919, 1011122811, -1136386606, -1136386606, -1221030748, -1215390919, -1249495107, 1011128180, -1125189627, -1214841163, -1084926640, 1063047003, -1214841163, -1136386606, -1223229771, -1203154020, -1156726498, -1198476264, -1212642140, 1013578459, -1136386606, -1127997998, -1084926640, 1063159478, -1136386606, 1062958654, -1084926640, -1136386606, 1040747617, -1217732213, -1115125579, 1040747214, -1115125579, -1223229771, 1022376699, -1199438337, -1249495107, -1125171910, -1200405241, -1217732213, -1197376753, 1013488265, 944604505, -1215390919, -1156705023, -1115125579, -1115125579, 919163804, -1207277189, 1051372795, 897988541, 921362827, -1125171910, -1214841163, 1063047574, -1214841163, -1084926640, 1024661085, -1136386606, -1127997998, 1040747617, -1115125579, -1217732213, 1040747080, -1115125579, -1228319844, -1115125579, -1115125579, 1051372795, -1214841163, -1217732213, 1011132475, -1215390919, -1241106499, -1218831725, -1249495107, 1003988334, -1143533969, -1232717891, -1215390919, -1143533969, 1062667620, -1217732213, -1084926640, -1136386606, -1228319844, -1230518868, -1217732213, 1011123885, -1115125579, 1040748556, -1115125579, -1208793849, -1115125579, 1040747818, -1115125579, -1214841163, -1102263091, -1115125579, -1115125579, 1051373433, -1210443117, 930850946, -1210443117, -1127997998, -1208793849, 953955186, 1020256596, -1190293815, -1162877428, -1206452555, -1232717891, -1192703828, 1016100142, -1192703828, -1131504302, -1127997998, -1214841163, -1190087656, -1163796551, -1193528462, 1020307599, -1206452555, -1206452555, -1131504302, -1206452555, 1054754948, -1093315231, -1084926640, -1093315231, 1067754119, -1136386606, -1127997998, 1019485650, -1136386606, -1136386606, 1040747617, -1115125579, -1217732213, 1040747214, -1115125579, -1223229771, 1022179131, -1249495107, -1199300898, -1199580608, -1125371626, -1115125579, -1115125579, 919163804, 1051372795, -1207826945, 916964780, 897988541, -1136386606, -1217732213, -1196826997, 944604505, 1013467864, -1156799512, -1215390919, -1136386606, -1223229771, -1202329387, -1198888581, -1157074390, 1013489338, -1213741652, -1223229771, -1202604265, -1156997081, -1198888581, -1213741652, -1136386606, 1013508666, -1084926640, -1125371626, -1214841163, -1214841163, 1063041332, -1084926640, -1093315231, -1136386606, -1084926640, 1074192179, -1136386606, -1218831725, -1207277189, -1236708452, -1249495107, -1249495107, -1127997998, 1019512493, -1224329283, -1212642140, -1167984681, -1173344800, 970698042, -1136386606, 1012196553, -1115125579, 1040747214, -1223229771, -1115125579, -1115125579, -1115125579, -1115125579, -1102263091, -1136386606, -1115125579, -1115125579, -1102263091, -1127997998, -1115125579, 1075742390, -1115125579, -1102263091, -1127997998, -1115125579, -1115125579, -1102263091, -1127997998, -1115125579, -1115125579, -1102263091, -1127997998, -1115125579, -1115125579, -1102263091, -1127997998, -1115125579, 1065353216, -1136386606, -1102263091, 1097859629, -1174306873, -1214841163, -1214841163, -1249495107, -1174289693, 992535267, -1165806595, -1165840955, -1196552119, -1217732213, -1136386606, -1215940675, -1163117946, 1011977510, 960488368, 968017983, -1136386606, -1223229771, -1212642140, -1167280306, 971660115, 1012239503, -1172880943, -1115125579, -1102263091, -1115125579, 906377149, 957189833, -1183490586, -1184246501, 1051382929};
localparam integer A_BRAMInd[0:664] = '{0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 5, 6, 1, 2, 3, 4, 5, 6, 0, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 3, 4, 5, 6, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 1, 3, 4, 5, 6, 7, 1, 2, 3, 4, 6, 0, 2, 3, 4, 5, 6, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 5, 6, 0, 3, 4, 5, 0, 1, 3, 4, 5, 6, 2, 3, 4, 5, 6, 7, 1, 3, 5, 0, 2, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 6, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 3, 4, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 3, 5, 6, 7, 0, 1, 2, 5, 1, 2, 4, 5, 7, 3, 4, 7, 2, 5, 7, 1, 2, 3, 4, 5, 7, 4, 7, 0, 1, 2, 3, 5, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 7, 0, 1, 2, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0};
localparam integer A_BRAMAddr[0:664] = '{0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 42, 42, 43, 43, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 48, 48, 48, 48, 49, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 51, 51, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 53, 53, 53, 53, 53, 53, 53, 53, 54, 54, 54, 54, 54, 54, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 57, 57, 57, 57, 58, 58, 58, 58, 58, 58, 59, 59, 59, 59, 59, 59, 60, 60, 60, 61, 61, 61, 61, 62, 62, 62, 62, 62, 62, 62, 62, 63, 63, 63, 63, 63, 63, 63, 63, 64, 64, 64, 64, 64, 64, 64, 64, 65, 65, 65, 65, 65, 65, 65, 66, 66, 66, 66, 66, 66, 66, 66, 67, 67, 67, 67, 67, 68, 68, 68, 68, 68, 68, 68, 69, 69, 69, 69, 69, 69, 69, 69, 70, 70, 70, 70, 71, 71, 71, 71, 71, 71, 71, 71, 72, 72, 72, 72, 72, 72, 72, 72, 73, 73, 73, 73, 73, 73, 73, 73, 74, 74, 74, 74, 74, 74, 74, 75, 75, 75, 75, 75, 75, 75, 76, 76, 76, 76, 76, 76, 77, 77, 77, 77, 77, 77, 77, 77, 78, 78, 78, 78, 78, 78, 78, 78, 79, 79, 79, 79, 79, 79, 79, 79, 80, 80, 80, 80, 80, 80, 80, 81, 81, 81, 81, 81, 81, 82, 82, 82, 82, 83, 83, 83, 83, 83, 84, 84, 84, 85, 85, 85, 86, 86, 86, 86, 86, 86, 87, 87, 88, 88, 88, 88, 88, 88, 89, 89, 89, 89, 89, 89, 89, 90, 90, 90, 90, 90, 90, 90, 90, 91, 91, 91, 91, 92, 92, 92, 92, 92, 93, 93, 94, 94, 94, 94, 96, 96, 96, 96, 96, 96, 96, 97, 97, 97, 97, 97, 97, 97, 97, 98, 98, 98, 98, 98, 98, 98, 99, 99, 99, 99, 99, 100, 100, 100, 100, 100, 100, 100, 100, 101};

//Conatant array to load the instruction BRAM
localparam integer total_instructions = 567;
localparam integer sub_instructions = 12;
localparam integer Inst[0:566][0:11] = '{{0, 0, 0, 0, 0, 0, 553648128, 540672, -2080374256, 2162688, 939526368, 2},{0, 0, -1818755072, 10764692, 0, 0, 595591300, 581896, 568, 2326528, 939524096, 2},{0, 0, 1151336448, 21518956, 0, 272629760, 394264670, 0, 1577058304, 1540096, 1883376064, 2},{0, 0, -1550319616, 10201366, 0, 0, 24, 889192448, -1710407304, 2523888, 416, 0},{0, 0, 1655439360, 18334126, 0, 272629760, 645922940, 630784, 0, 134217728, -130742623, 1},{0, 0, 1244397568, 12309066, 0, 0, 109170688, 106612, 0, 2556896, 1879050176, 2},{0, 0, -1827667968, 22656340, 0, 125829120, 251658264, 402653184, 805306984, 427216, 0, 0},{0, 0, -1557397504, 18301367, 0, 0, 343933052, 335872, 974356480, 950272, 1879050208, 2},{0, 0, 1655439360, 21576974, 0, 121634816, 251658288, 237568, 2080374784, 0, -937490496, 0},{0, 0, -1842610176, 15017623, 0, 318767104, 82, 335872, 0, -1945140688, 1744831456, 2},{0, 0, -1827405824, 14000886, 0, 260046848, 154, 196916, 805912872, 2064384, 0, 0},{0, 0, -1667497984, 17281782, 0, 260046848, 394264660, 0, 1141883152, 0, -2144665600, 1},{0, 0, -1306001408, 16499145, 0, 0, 84, 434344, 1778893136, -1409286144, 992, 0},{0, 0, 1419509760, 20459215, 0, 0, 0, 1308926200, 1242137072, 1245184, 1879048192, 2},{0, 0, -2070151168, 18103699, 0, 0, 67264528, 73880, 1174405192, 0, 1120, 0},{0, 0, 1419771904, 22665870, 0, 0, 562036888, 637812736, 1140850936, 874611296, 407110625, 2},{393216, 114768, 1419509776, 1393995472, 1548810401, 539408, 557981764, 1242104104, -2062417388, 539231056, 1077217521, 2},{470024512, 100663296, 0, -412437216, 1739362953, 327891728, 600068229, 1174991000, 301990272, 2343680, 2015822112, 2},{384, 114688, 16404, 15017568, 1222420480, 223165482, 461410399, 201719856, 1594638408, -1005060096, 339085776, 2},{-2147483648, 98370, 28, 825808384, 1496100769, 102179416, 528765088, 797434176, -1694170708, 1680146752, 1476395440, 2},{327680, -1073741824, 28688, 1828105952, 1278249113, 38944042, 650440862, 151519548, -1710964584, -702545408, -61863856, 1},{274432, 87556096, 0, 829997536, 1498737001, 1275288, 247519232, 537509988, 838877296, 69158120, 1879116256, 0},{-2147483264, 117440578, 0, -1326142176, 1429771145, 264780836, 662700093, 1300750412, 637534404, 1074184672, -265681599, 0},{262144, 84992, 28, 1463222272, 2074380961, 134755172, 348389438, 254032, -1660460984, 2014315520, 1343555568, 0},{384, 65536, 21376, 714711552, 1529927529, 734756, 360845371, 587473036, 2098119128, 1410336, -65436576, 0},{384, 70778880, 20480, 557139264, 2058664057, 155989284, 209866835, 84402180, 838942728, 336708088, 1816134880, 2},{469762432, 83886144, -2147483648, 821413235, 1271441745, 202259754, 293855387, 1040388348, 1610613036, 2080768, 536872321, 1},{0, 65616, -2013240448, 385135925, 1411963033, 97402344, 192938090, 486891652, 2131427604, 604930192, 1546683776, 1},{283115520, 98304, 1610612756, -1317390991, 1546170265, 349584932, 310411420, 348374, 1058259104, -1607892672, 1074333040, 1},{417333248, 81984, 0, 788965024, 1201711969, 43269676, 302161990, 705155222, 1292010100, -1878687728, 671154496, 1},{470024512, 98304, 0, -1865099744, 1708960929, 4860908, 323100689, 16855168, 1191821944, 1310800, 1076035744, 1},{469762048, 67, -1476394988, 427341129, 1815910465, 51392038, 553865354, 528765164, -1308622540, 203261328, 806160817, 2},{136, 83902464, 12288, 647739808, 1079294049, 146186775, 335712391, 0, -2030042824, -1541750096, 608700640, 2},{140509184, 18432, 20480, 1462272000, -1606371167, 277720594, 92344458, 1493766442, -1862115248, 329104, 1007747072, 1},{268763136, 0, 8192, 722894848, 1481685065, 1488984, 79908996, 419532884, 704643460, 201326592, 2082080417, 2},{67109056, 34816, 20, 637534208, -1606112911, 767530, 595918959, 1241911336, 1661280760, 941555872, 817, 0},{67109120, 80, 0, 637534208, 1096115049, 9461795, 662700051, 1074319372, 156, 98304, -134215232, 1},{0, 51200, 8212, 649363456, -2133021511, 55857186, 159432860, 201588788, 1090543816, 2556400, -2078736336, 2},{268435456, 0, 0, 827907680, -1857444959, 160850016, 243310636, 1057124504, 2081063028, 328048, 960, 0},{0, 1610612736, 17032, 460962880, -525290063, 84582434, 302071878, 507984, -2146893824, 1108476496, -1408596655, 0},{268435524, 80, 0, 460969568, 1448644513, 137269484, 58720319, 721711272, 1023410460, 201392128, 403112000, 0},{-1744764928, 34866, 0, 1744830464, 1713425225, 1153044, 281428162, 92287368, -1526636068, -1876623360, 675415233, 3},{12352, 53018624, 8192, 278953984, 1236055385, 197938732, 214165579, 805626004, 17563792, -1676427256, 69075520, 2},{8, 36175968, 4108, 1610612736, 2024069201, 99327135, 335700065, 755318784, 704872684, 873873560, 604899344, 1},{70, 32832, 20480, 805306368, 740650865, 141864483, 109072471, 722059284, 1494433956, 404439312, 1280246304, 0},{327872, 67125248, 8, 12179040, -188434432, 697188, 356659367, 73864, -1627389664, 738246816, 872416528, 1},{256, 83886080, 24576, -948404224, 816726660, 416124971, 33558531, 16809984, -972308328, 1409467152, 476055072, 1},{131072, 1654784, 4608, 1901646400, -155666615, 323716628, 331362398, 839270720, -1290747368, 1143489160, 202211457, 1},{209715200, 16809984, 0, 15777824, 1767148032, 80984803, 159383696, 319254530, 1829896768, 606192752, 877201633, 2},{128, 16777280, 12, 15777824, -707180288, 127176172, 260157519, 402907244, 1460044492, 673464736, 1209599280, 0},{196608, 0, 8192, 33554432, 399176794, 248728923, 147038290, 486694912, 1812415028, 1411482464, 1680475840, 0},{0, 0, 193073408, -2046416851, -64563108, 1412586, 671412404, 729376, -1575746960, -1875770240, -1273329663, 1},{201326720, 0, 4112, 423012352, 122197593, 269845481, 532734113, 1090605056, 512, 67568624, 1544618001, 2},{73662474, 33554432, 0, 805306368, 1522644809, 57371736, 104960159, 84414478, 1511424720, -66994096, -802289632, 0},{67240192, 81920, 12288, 1397792800, -668370831, 93294110, 272887885, 436416608, 1426555120, 1544355840, -1539307024, 0},{141568, 1572864, 67108864, 10127023, 1549568768, 135044206, 88164393, 537166084, 2113929728, 68108664, 404686817, 1},{0, 16809984, 0, 100663296, -1681833838, 59471074, 461373442, 352468, 1224785920, 873612160, 1476592096, 1},{196608, -2130706432, 8, -1621622784, -1253506995, 106208110, 63234202, 1325604864, -939523384, -1711192848, -2142437264, 2},{67239936, 0, 0, 24707072, -1808137472, 148222818, 843251808, 84693184, -1795079496, 1477378608, 540608161, 1},{-2147483648, 17, 144179200, 1362154550, 405100731, 21724695, 109076554, 310702100, 201326980, 458848, 1076232448, 0},{67315712, 0, 16, 729392832, 1461758569, 59547802, 180377681, 373120, 1443529104, -2079883056, -1741684527, 1},{256, 0, 4096, 12156928, -700849664, 143673902, 84127745, 294952, 68075800, 67683344, 2084503617, 2},{272384, 33554432, 4, 489705472, -1765088431, 1017174, 12601478, 557076, 352322080, 376832, 805700752, 2},{128, 575568, 0, 1889107968, 1545640001, 307242156, 612671687, 352919848, -1055858148, 705304, -1476395008, 0},{67108864, 1073807440, 0, 1845493760, 1246533009, 160515620, 327155846, 654725496, -1861172668, 305071216, -1606153680, 0},{0, 0, 8196, 8388608, 2052712704, 281832675, 150994983, 906412080, -2013101536, -2147483648, 1279592752, 2},{268439552, 100683264, 20, 1689325024, 1195411849, 1351214, 230815816, 570978596, 890085664, -1474608208, 1344472784, 2},{209715264, 0, 20, 2457600, 1144332288, 1084838, 746864757, 1124249890, -1878474208, 603979776, 1211762705, 2},{0, 50332160, 0, -1006632960, -440257115, 382303760, 226885686, 196992, -1592500224, 1681016256, -665058464, 0},{73862, 0, 20480, -245792768, 1264471370, 73933480, 121739393, 1393172728, 524, 2720992, -732821056, 0},{-2147483328, 35859, 12800, 0, 884037632, 130837605, 801239167, 511926628, -2096651564, 1680867328, 1950385024, 1},{0, 0, 4104, 24805376, -1258291200, 18049828, 25530494, 17301520, 1074233556, 1744961536, -1140718863, 0},{262144, 50331648, 0, 379117152, 1632668841, 227440741, 4305006, 536680, 872415664, 1229664, -536870912, 0},{131328, 49152, 4, 268435456, 1238999209, 328232412, 365031475, 822730948, 118719080, 1605632, 496, 1},{283443584, 0, 8192, -1500872704, -265244319, 26378350, 406863969, 397434, 1208074696, -669908128, 738198656, 3},{256, 16, 402666120, 10596462, -1140215808, 232238020, 725671947, 234995904, 1645052604, -669483008, 606504752, 1},{0, -2147483136, 12713992, 17844245, -1137545728, 39288366, 92274784, 503726152, 486646024, -2046230336, 1344405777, 0},{268763136, 16777216, 8192, 436207616, 1613951906, 1084005, 88182822, 436293656, 268861496, 1342685280, 1678246112, 1},{0, 16826368, 8704, 482017280, 1235783753, 206548058, 499318932, 1577664632, 84410944, 471909856, 738625089, 1},{0, 1124073472, 4, 738197504, 1012837012, 875615, 654626882, 554209568, -1845001664, 438518928, 1213139089, 2},{69638, 0, 16384, 436207616, 1419931204, 309427625, 616867883, 549124, 560, 2229264, -1538914175, 0},{65536, 80, 8208, 10563648, 671088640, 244145363, 331571326, 504090624, 303054932, 1210089472, 605226000, 2},{201326592, 67125248, 8192, 22118400, 473091840, 244019823, 302120997, 446584, -1995964176, 1393200, 740361216, 2},{0, 0, 4096, -1006632960, 80847036, 1398303, 402653284, 1661755592, -1039072696, 3180064, 1413745728, 2},{139456, 0, 4, 620019744, 1193840009, 106145176, 575015093, 245760, 905969928, 1917360, -669382352, 0},{64, 33554480, 0, 0, 1990274560, 340825617, 679477303, 606496, 740, -64076848, 1480524656, 2},{256, 32768, 0, 805306368, 877748585, 13913573, 226492479, 67125608, -1493138788, -2144534496, -805306303, 0},{320, 0, 16384, 1727431008, 1230803297, 206848084, 361041929, 262336, 1040891904, 1377264, 338823744, 0},{65536, 33554432, 12, -2147483648, -899782253, 1403550, 541393024, 442624, -1676836432, 1140999120, 3607377, 2},{67108864, 33554432, 12800, 805896192, -439544215, 202406506, 301989986, 217324, 1980285208, 1852192, -467630944, 0},{201326592, 19496992, 16, 0, 89844992, 949481, 125829150, 405564, 1224982924, 1009238600, -2079325040, 2},{335951872, 16777250, 0, -1509949440, 1263577433, 386608104, 121661556, 243388612, 252150220, 1884720, -802158784, 1},{0, 1024, 4096, 19988480, -64902656, 1527340, 671133718, 235151396, 1896636664, 492768, -1001324064, 1},{134217728, 50331648, 4112, 0, -727044972, 160800168, 335679540, 235032680, 202129800, -2147073776, -1675033968, 1},{0, 49153, 6029312, 17288214, 1958098944, 1400361, 125886542, 126410908, 286752980, 1278208, 805307584, 1},{192, 1073741824, 4, -2147483648, -1422847108, 286567256, 411213973, 755531776, -1643363832, -903379952, 3015728, 2},{0, 52985856, 134221840, 21475374, -2008500480, 85043802, 419516483, 409792, -1828716376, -534461368, 2084046992, 2},{262144, 16, 0, 0, 975473408, 1097061, 457457684, 536848, 369099316, 336135248, 1342769281, 0},{0, 32768, 4, 0, -1496492702, 404114326, 629276752, 328064, -2095922648, 335544320, 2492273, 1},{134, 65616, 0, 58294272, 1211937962, 250760598, 520187977, 1493844292, -1994866100, 269534304, 538446017, 3},{201326592, 33570816, 0, 10125312, 1227451648, 55544359, 101, 815376, -1022295504, 405882000, 677054753, 2},{0, 16809984, 0, 13959168, -129112064, 638486, 511959166, 587202560, 923795920, -2146581552, 138019920, 2},{0, 83937280, 4096, -402653184, 1409466986, 625695, 612761763, 1678540800, 2063639112, 674250784, 1548683745, 2},{201326592, 32, 0, 10782112, 92274688, 181513385, 268656702, 741556, 1846231076, -602176864, 1610613648, 1},{65792, 0, 8192, 493920288, 1448264537, 5205207, 365166701, 442424, -1978269696, 337772816, -1806169519, 1},{0, 48, 4, 2785856, 1009618432, 227130331, 385876040, 990232576, 492, -1877867648, -1071314384, 1},{0, 33554432, 0, -1052180480, 1993965962, 131488337, 427954242, 475276, -1844346472, 404309056, -805304031, 1},{209715264, 0, 8192, 686096384, 2066591617, 227056811, 620863519, 956428486, 520520264, 1867776, -2078668448, 0},{0, 0, 4104, 0, -1697510912, 114080862, 276869138, 855761100, -1157382024, 806223872, -601880752, 1},{350224396, 33554496, 268439552, -1729019822, 1238813625, 112478434, 453361687, 788746266, 1912930700, 1946665872, -1944714559, 2},{0, 32768, 4096, 0, -180974080, 1411794, 102, 1208360960, 588022168, 1131296, 1278345216, 1},{134479936, 2719792, 0, 1879048192, 1203803676, 340366162, 415526991, 822407168, -1625849100, 1208501496, -1874852287, 1},{128, 16, 0, 0, -1784534528, 332377646, 411041929, 319572, 1309245964, 1076330832, 1947469409, 1},{2048, 0, 8, 335544320, -111310067, 332221660, 180562056, 65536, -1609317624, 402949648, 1476921104, 0},{131328, 16777216, 12288, 560005120, -148799383, 336157870, 574824641, 401408, -1575763968, 2278640, -1674376672, 0},{131072, 16, 12800, 0, 618506752, 89619371, 633671761, 1258504192, -1777352148, 1343062352, 202933088, 1},{0, 35651584, 0, -1040187392, 641241515, 114122197, 570630244, 213152, 392, -1742519144, 605816096, 3},{0, 16, 0, 2752512, 618010112, 366172847, 176, 1074491776, 2113946164, -1877867616, 134219584, 3},{335740928, 0, 8208, -326533120, -525762373, 306862946, 516198600, 20656, -938065128, -2078931824, -1805383183, 2},{256, 0, 20484, -335544320, -609176717, 349198954, 87, 823524, -1508655104, -2078637552, 1681459536, 1},{136, 16777216, 268455936, 3189837, -914358272, 271482322, 151044161, 373068, -1508670824, 1819952, -1139602976, 1},{262144, 1040, 0, 0, -105295872, 332704346, 390373524, 923197440, -1324261236, -601586832, -2143876640, 2},{201326592, 16842752, 0, 19302400, -1537894912, 181095534, 377729184, 487604, -1828126248, 1008484928, 743507777, 1},{196672, 32768, 0, -1073741824, 2052680019, 63991143, 432078915, 131088, -1929117568, 0, 671089152, 0},{-1744764928, 65538, 8, -1433829376, 1211937401, 135735966, 222597142, 260173864, 521290188, 0, 1344342384, 2},{67108864, 50331648, 0, 10190848, 822083584, 1407533, 218173466, 436629804, -1777188704, 934240, 336986656, 1},{0, 536903680, 0, 21528576, 112849664, 46839123, 620793886, 302112768, 1930575952, 1510474016, 1477184432, 2},{196736, 16384, 0, -805306368, 81415331, 269331567, 792744039, 1091108864, 1695564528, 1654896, -1879047968, 2},{0, 0, 8, -2147483648, 2023940484, 63613791, 318849110, 352321536, 1476641080, 1441792, -2147482032, 0},{256, 1610612736, 8, 1073741824, 1732411789, 22510105, 234897545, 1510178920, -1039269840, -838662752, -1070134768, 1},{0, 17408, 0, 1580662784, 2018145346, 47033433, 83886098, 69812, -1593647016, 739836096, 1881933376, 1},{0, 0, 4104, 12910592, -1808871424, 286761830, 17141922, 0, -1559150592, 2261040, -1671820751, 1},{0, 16777248, 16384, -973078528, 649260978, 248877673, 43, 1644961932, 1678688860, -938621424, 738200640, 2},{128, 0, 4608, 15040512, 1227395328, 286236122, 101, 524324, -1945862144, 2294048, -463370959, 0},{192, 32, 0, 0, 2001297664, 891865, 177, 1678213120, 2046820820, 1916928, -664729280, 1},{134217792, 100728832, 20, 1184923648, 1815656586, 1189392, 16777363, 50696192, 1863156264, -468663216, 608502832, 3},{0, 0, 0, 0, -1741823744, 1358938, 167, 491520, -1509015552, 2588672, -402651392, 1},{268435456, 32, 20, 268435456, 1279039633, 942164, 0, 252112964, -1610333540, 1076364144, -1677720399, 0},{128, 0, 135925760, 11579438, 0, 26184896, 149, 483356, 1845494320, -534576256, -2075851616, 2},{201392128, 0, 8704, 637534208, -1740029767, 403403608, 382087234, 1661423616, 570671240, -2079260144, -1945795520, 2},{134414336, 16, 16384, -536870912, -698783117, 118603116, 138449042, 135280, 369213572, 738361344, 201785872, 1},{262144, 0, 4, 720896, 1464637184, 615383, 222355522, 973078528, 1913504200, -1811381344, 270598544, 1},{134217728, 16777216, 0, 1073741824, -128374683, 114121820, 218103880, 618496, 1208959464, 1879786064, -668924064, 1},{0, 33554432, 4480, -1711276032, -1742656845, 1549022, 545366190, 1577828352, 907149460, 67650944, 1682670432, 0},{192, 16, 8, 21004288, -114643456, 165043042, 327405757, 738287616, 2046968332, 1073988112, 1476397648, 0},{140509184, 16448, 96731136, 21054507, -629145600, 13139100, 754978868, 453308502, 1493271308, 271417552, -2080373920, 0},{131072, 67158016, 0, 1540096, -701837056, 1551080, 239165622, 402735280, 1896547028, 1654960, -1206645888, 0},{0, 0, 4096, 20414464, -1808383488, 89557674, 8474802, 565332, 33554432, 67519776, 1946356128, 1},{0, 34816, 268435456, -1048979854, -1582923342, 1472026, 427909220, 417792, -1962106880, 1343816048, -667745248, 1},{67108864, 32, 0, -2147483648, -900101822, 215309156, 537247844, 1443639500, 1678492436, 1476919376, -2141387167, 0},{0, 512, 16, -1799091584, -187836493, 30108778, 33579060, 229408, 621912128, 537133056, -402323120, 0},{134217920, 0, 4096, -1879048192, 1507757205, 9915415, 507818185, 504196, -1978121640, 1867792, -466155200, 1},{0, 0, 0, 20415936, -1856135168, 1070424, 0, 0, -1543503208, 0, -2013265920, 2},{-2147352576, 83984403, 12304, -1342177280, 1279295601, 4730396, 482385926, 931282984, -1593540156, 2637888, -334296560, 1},{0, 0, 0, 0, 1421767168, 349616991, 148, 1392652512, 169083328, 673710080, 939526497, 0},{131072, 16, 0, -2030023680, -866555325, 1146338, 499122182, 1628200964, -1575747020, 1075593216, -2013001183, 2},{0, 16777264, 16392, 1073741824, -148804972, 1481296, 10, 167772160, 140, 470892720, 1409287248, 2},{128, 0, 0, 0, 1610612736, 311265367, 57, 922870060, 571343448, -535756800, 1481245760, 2},{-2147483648, 0, 8192, -2036256704, -1713559436, 17533920, 41943054, 965386240, -1409154604, 2786656, 337971776, 1},{262144, 1073741840, 0, 607420416, 1193842785, 408337371, 549634136, 1225441280, -1006632468, -299171840, 805307280, 0},{67371456, 32848, 24, 1879048192, -1990937076, 1534872, 331362383, 923521264, 922812772, 741097472, 1342177808, 0},{65536, 64, 0, 0, 472711168, 1424359, 516079694, 268566540, 1342619700, -1609728000, 402784768, 0},{268435456, 16777216, 0, 821430656, 1732596393, 543959, 327155792, 364544, -1945796000, 1479393280, 1613299856, 2},{402981120, 32, 4096, 503316480, 1814089817, 1483356, 180539435, 738767024, -1543471012, 203948032, -1137833072, 0},{0, 0, 12288, -1006632960, 473530715, 89496171, 327155903, 285351936, 1207960024, 1075413632, -736688896, 2},{65536, 67108864, 8832, -1061093376, 1187103565, 198270101, 432099512, 167772160, 603979920, 541024, -1673428288, 1},{128, 0, 12, 0, 1457185024, 21924885, 134602855, 269205504, 692, 525456, 1611138672, 2},{-2071986176, 2, 12288, -1006632960, -903825331, 164785506, 16777296, 1166086534, 100663364, -1543503872, -332200352, 0},{67108864, 32, 0, 10780672, 1971322880, 18131885, 633425932, 117911812, -2113929188, 0, 135725792, 2},{134414336, 16, 0, 0, 1429803776, 395754579, 692306088, 956985720, -1845493100, 2670592, 0, 0},{144703488, 64, 4096, 805306368, 1549056177, 1275362, 754974730, 1442992354, 452, 872564064, -1677718688, 0},{201392128, 0, 8, 0, -1258291200, 365802600, 700448935, 1157689344, -1946156496, 1879080960, -535230095, 2},{196608, 16384, 8, 0, -1782960128, 1533456, 834670592, 923213828, -1559347152, 1610843520, 609749553, 0},{0, 83886080, 16, 33554432, 901657188, 633683, 478396616, 940343684, 385909192, 269566848, -402389936, 1},{67305472, 67108864, 8192, 1745256448, -170514300, 1219986, 147050664, 1024028896, 369098840, 1229344, 1547437920, 2},{128, 512, 0, 17235968, -723885312, 403795284, 142606501, 67125248, 286630024, -2012741632, 536872353, 0},{67108992, 0, 12288, 10551296, -902897664, 4756576, 83886169, 34263284, 488, 134578176, -67107776, 2},{64, 2128, 0, 0, -1447919104, 185318496, 121, 1677738216, 151445724, -2078473648, 671088737, 3},{134217728, 16384, 0, 3899392, -643153920, 1137176, 234881080, 135168, 1359397080, 917504, -534969472, 0},{65536, 49184, 0, -738197504, -81654717, 408191592, 591605792, 50462744, 755106404, 0, 1281491200, 1},{134217792, 52428800, 0, 23676000, 936679424, 404183637, 838860891, 1678397440, 1342177600, -2013150408, 1946158944, 1},{0, 18350080, 0, 14729248, -1325400064, 1162516, 402681856, 143688, 738197680, 403980664, -1874788128, 2},{0, 16777216, 8192, 14729248, -1718970368, 679248, 436207616, 872546696, 148, -2079636688, -335541183, 2},{0, -2097152000, 8, 1638400, -633038848, 415915234, 792723552, 704536, -1172995304, -838582272, -396293744, 2},{0, 0, 4, 0, 958582272, 370167263, 427819110, 1644216708, 117441032, -872184288, -1073609424, 2},{0, 0, 4, -2144862208, -1680771484, 374185040, 788529332, 393572, 768, 1946189824, 1348272881, 2},{64, 1610612736, 8, 0, -886682718, 1274926, 109052019, 0, -1409286096, 1442840576, -671086671, 2},{0, 0, 0, 0, 0, 565341, 587587634, 573440, 48, 671350784, -134217471, 2},{0, 1, 4, 18960448, 101111808, 60119573, 813695144, 1182851072, 67109572, -2077196288, 2014120849, 0},{134217728, 51200, 4, -2128510976, -1168599029, 1526296, 209715200, 471040, 252584672, 1882062848, -805303535, 0},{196608, 64, 8196, 0, 1174405120, 189482007, 482345161, 956768256, 1879048284, 0, -335544176, 1},{134217728, 0, 4112, 0, 1275068416, 1143982, 516145272, 185249792, 1879048968, 808517632, -468974160, 1},{65536, 0, 0, 0, 363987456, 1406355, 147030016, 1459617792, 369098788, 939591008, 1879900352, 0},{67108864, 0, 16384, 2556288, -1462462464, 543450, 0, 185053256, 144, 98304, 1811939328, 1},{67108864, 0, 0, 2490368, 0, 1084608, 0, 479300, 939524096, 0, 738197504, 3},{72, 80, 12, 2209888, 0, 70460928, 57, 0, 28, -805306368, -332856432, 0},{0, 18512, 256, 0, 1275068416, 601622, 0, 1627873680, 285876548, -267223040, 338985696, 3},{0, 65616, 0, 1073741824, 1546426524, 1204308, 50331680, 1409982464, 755630260, 229376, 1207960864, 1},{67371008, 33554432, 0, 0, -180053915, 1160336, 138412122, 675840, 738197824, 1546568048, 1881998976, 1},{4194304, 0, 0, 0, -1809186560, 750444, 0, 51138770, 134217904, 271220736, -402651264, 1},{75497472, 32768, 0, 0, 70293504, 756629, 199, 708870, -1157513216, 0, -1610612736, 1},{68, 0, 0, 8457696, 0, 216006656, 411041969, 51003652, 788, 0, -805303744, 2},{192, 0, 8, 0, 1277305088, 695429, 142672061, 114756, -1811938556, 805306368, 2993, 0},{268763136, 16, 0, -1342177280, 1546426372, 1289500, 591396864, 822661316, -1174404428, 1949204480, 2929, 0},{268435456, 16809984, 0, 0, 369098752, 760727, 587259904, 234942828, -1189592480, 1812219312, -67106431, 2},{0, 50331648, 256, 1540096, 380276736, 369863895, 218103860, 16412, 64, 2900096, 2085980928, 0},{0, 16777216, 0, -1342177280, 730234893, 891925, 469762048, 50905088, -1811938624, 3032448, 1476396448, 2},{0, 0, 4, 0, 609304576, 887837, 721420288, 1443053596, 404161296, 3014656, 1488, 0},{268435456, 32848, 4, 14729280, 662700032, 1154329, 50331769, 94208, -988446700, 0, 400, 0},{268435584, 0, 0, 0, 0, 118464576, 113, 28716, 2013266064, 393216, 1611858384, 0},{0, 67190784, 0, 805306368, 912046193, 1088081, 190, 67260428, 956350480, 269369408, 542769248, 0},{0, 0, 0, 503316480, 950144340, 415866263, 56, 811396, -1342177264, 917504, -1810035968, 0},{0, 16777216, 0, 0, 123308288, 1220053, 0, 1493172224, 1392509696, 1720320, 0, 3},{196608, 33570816, 0, 0, 0, 560128, 843055223, 0, 789200896, 1983120, 0, 0},{4390912, 0, 4, 15774752, 0, 0, 62914560, 700754, 771751936, -1207959552, 1328, 0},{131072, 0, 4096, 11581440, 0, 0, 440401920, 0, 2013724672, 770048, 1946157056, 1},{0, 1104, 16384, 0, 0, 948288, 0, 0, 152395836, 0, -1543503872, 1},{0, 0, 0, 0, 0, 0, 436236288, 1443266904, 235012152, 2949248, 674496512, 0},{0, 16, 0, 89587712, 130626658, 1148123, 34, 675840, 748, 0, -1879048192, 0},{0, 17874944, 0, 23076864, 0, 0, 146800640, 118177792, -1224736048, 2475208, 0, 0},{262144, 16777216, 0, 0, 0, 1084544, 817889280, 122880, -1157627784, 3063808, 0, 0},{0, 16777248, 0, 0, 536870912, 99843, 813694976, 24972, 612, 2999680, 536870912, 3},{201326592, 1, 0, 0, 545259520, 1286683, 0, 1552650312, -1241268156, 2459056, 2400, 0},{-2013265920, 65538, 4096, 10530848, 1275068416, 883622, 813694976, 1653027216, 420954820, 3048224, 1550123008, 2},{0, 16384, 0, 0, -679477248, 1286744, 726011904, 802816, -1190362392, 3048992, 0, 0},{0, 0, 0, 0, -134217728, 896152, 838861000, 1644863488, -1476197700, 0, 384, 0},{0, 48, 8, 1376256, -117440512, 1346972, 0, 1543503872, -1207516700, 98304, -1677720656, 0},{0, 33554448, 0, 3538944, 0, 949312, 830472383, 1644167168, 36, 147456, 928, 0},{0, 16384, 8192, 10551296, 0, 1345536, 0, 0, -1324646400, 1508160, -335541248, 0},{0, 83951616, 0, 327680, 1546694400, 796186, 0, 453173616, 1394016624, 1359872, 0, 0},{0, 81920, 16, 0, 1547737088, 1019108, 0, 0, 788529152, 0, 1488, 0},{0, 0, 0, 0, 0, 0, 112, 466944, 771751936, 1966080, 1472, 0},{0, 0, 0, 0, -536870912, 1463448, 0, 0, 0, 0, 0, 0},{262144, 0, 0, 0, 0, 0, 62914560, 688128, 1375731776, 1703936, 0, 0},{200, 16384, 20480, 16809984, 1275068416, 74215588, 58720437, 1443549216, 285213368, 262144, -1811939328, 0},{0, 0, 0, 0, 1233125376, 72459289, 796946468, 0, 720, 0, -1744830464, 0},{0, 0, 0, 0, 1946157056, 1092909, 180, 741376, -1274986496, 0, 0, 0},{67108864, 0, 0, 0, 0, 395214208, 150, 749868, -1744829732, 2490368, 0, 0},{64, 83886080, 16, 0, 1197258752, 76754328, 177, 0, 0, 2473984, 605161840, 3},{0, 0, 0, 0, 0, 1525824, 629145788, 614400, -1224736768, 1671168, -134215328, 2},{0, 16384, 0, 0, -1442473984, 1462820, 0, 0, -1156021664, 2491568, 738197504, 3},{0, 67108880, 0, 491520, 0, 814080, 0, 1527415148, -1241513236, 409856, -1879047680, 0},{0, 65536, 0, 0, -1463222016, 945372, 201, 0, 117899264, 0, 0, 0},{0, 0, 16, 0, 0, 32256, 0, 1560281088, -1174404380, -872415232, 944, 0},{0, 64, 0, 0, 0, 941120, 199, 376832, 102105860, 1744962944, -805306239, 2},{0, 17408, 0, 589824, -408302592, 553690, 192937984, 376832, 1762370272, 917504, 0, 0},{0, 0, 0, 2688640, 0, 1073152, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 478150770, 0, 480, 0, 928, 0},{0, 0, 0, 20994048, 0, 1069120, 0, 471040, 0, 0, 0, 0},{0, 64, 0, 0, 0, 0, 104, 0, -1476394940, 393216, 0, 0},{0, 0, 0, 23068672, 0, 942144, 440754176, 704512, 268435520, 0, 0, 0},{0, 0, 0, 1507328, 0, 1213760, 0, 147456, 700, 393216, 0, 0},{0, 0, 0, 0, 0, 1204288, 801112064, 57344, 720, 0, 0, 0},{0, 0, 0, 0, 0, 1085440, 0, 0, 0, 0, 0, 0},{0, 16384, 8, 0, 0, 0, 151, 0, -1728053248, 0, 3056, 0},{0, 0, 0, 0, 0, 0, 150, 0, 0, 0, 624, 0},{142671872, 0, 0, 23101440, 0, 0, 633339904, 766346, 0, 0, -67108864, 2},{0, 0, 0, 0, 0, 0, 134623264, 802816, 612, 0, 536870912, 3},{134217728, 16, 0, 0, 1074190336, 1413635, 838860800, 700808, 732, 0, 671088640, 3},{0, 0, 0, 0, 0, 1350144, 0, 0, 0, 0, -201326592, 2},{256, 0, 0, 0, 0, 0, 93, 67108864, 134218476, 0, 0, 0},{0, -1577041920, 16384, 17905728, 0, 0, 0, 761856, -1325399320, 1644314624, 2083785552, 1},{0, 0, 0, 0, 0, 1068160, 0, 757760, 0, 0, 0, 0},{262464, 0, 0, 0, 0, 0, 482345075, 753664, 0, 0, -268434528, 2},{0, 0, 0, 0, 0, 240275968, 478150776, 696320, 0, 1409286144, -329971807, 1},{256, 0, 0, 0, 1171974656, 252296339, 478150761, 0, 0, 0, -402653184, 1},{268435456, 0, 0, 0, 0, 1548800, 708837480, 69632, 1946157520, 0, 0, 0},{0, 0, 0, 0, 0, 963584, 725614592, 704544, 696, 0, 608, 0},{0, 0, 0, 10485760, 0, 1219584, 796917760, 737312, 64, 0, -1677721600, 0},{0, 0, 0, 0, 0, 1219877, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{256, 0, 0, 0, 0, 0, 151, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 150, 0, -1744829856, 0, -134214688, 2},{0, 0, 0, 0, 1744830464, 570013, 34, 0, 0, 0, -1879048192, 0},{67108864, 0, 0, 0, -2130706432, 112130, 0, 749568, 0, 0, 603979776, 3},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 738197504, 3},{0, 81984, 0, 0, 0, 0, 0, 0, 150994980, 0, 0, 0},{0, 0, 0, 0, 0, 369098752, 104, 1476395008, -1342111712, 0, 0, 0},{0, 0, 0, 0, 193124352, 949341, 190, 765952, 32, 0, 2880, 0},{0, 0, 0, 0, 0, 689536, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -201326592, 2},{0, 1073741824, 4, 0, 0, 0, 0, 700416, 0, -167772160, 2736, 0},{0, 0, 0, 0, 0, 0, 0, 475136, 0, 0, -335544320, 1},{0, 0, 16, 18874368, 0, 0, 0, 0, 468, -201326592, -402652560, 1},{0, 0, 0, 11796480, 0, 0, 704643072, 696320, 134218428, 1275068416, 2880, 0},{0, 0, 0, 0, -528482304, 1334420, 801112064, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 637534208, 622592, 0, 0, 0, 0},{0, 16, 0, 18927648, 0, 0, 0, 0, 612, 1275068416, 3056, 0},{0, 0, 0, 0, 0, 22592, 767557632, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{131136, 0, 0, 0, 0, 0, 784335025, 0, 708, 0, 0, 0},{0, 0, 0, 0, 0, 0, 191, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 780140544, 0, 0, 0, 0, 0},{268435456, 0, 0, 0, 0, 1320448, 0, 479232, 0, 0, 0, 0},{0, 0, 16, 0, 0, 0, 494927990, 475136, 0, 0, 1968, 0},{0, 0, 0, 0, 0, 1348992, 754974720, 0, 0, -201326592, 1744833184, 0},{0, 0, 0, 0, -2139095040, 677928, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 172, 0, 640, 0, 3040, 0},{268763136, 0, 0, 0, 1277728768, 1060396, 641728512, 626688, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 637534380, 1460240384, 640, 1140850688, -268433503, 2},{0, 0, 0, 0, 631324672, 1483873, 797229056, 0, 0, 0, 3040, 0},{0, 0, 0, 0, 0, 699648, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 187, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -536870912, 1},{0, 0, 0, 8388608, 0, 0, 119, 0, 0, 0, 0, 0},{64, 0, 0, 0, 0, 0, 181, 700416, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 33554432, 4096, 0, 0, 0, 0, 0, 652, 3129344, -1140850688, 2},{0, 0, 0, 0, 0, 0, 0, 0, -1577057656, 2654208, 0, 0},{134217728, 0, 134217732, 12630064, 0, 0, 0, 782336, 700, 0, 2608, 0},{0, 0, 0, 0, 0, 0, 801112064, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 186, 0, 0, 0, 0, 0},{0, 0, 16384, 0, 0, 1451520, 0, 0, 0, 0, -469762048, 1},{0, 0, 0, 0, 0, 0, 511705088, 499712, 0, 0, -536870912, 1},{0, 0, 0, 0, 0, 1197312, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 679936, 656, 0, -1207959552, 2},{0, 67190880, 0, 1879048192, 1279842369, 1062416, 0, 0, -1560280436, 2670592, 0, 0},{0, 0, 0, 0, 0, 0, 688205990, 672076, -1577057648, 2654208, 0, 0},{0, 0, 0, 603979776, -893266813, 1275302, 796917760, 1358954496, -1577057608, 3114256, -1207959552, 2},{0, 0, 0, 1879048192, -333303709, 822552, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3024, 0},{0, 0, 0, 0, 0, 0, 122, 0, 0, 0, -268435456, 1},{0, 0, 0, 23076864, 0, 0, 515899392, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 1124073472, 4, 0, 0, 0, 0, 0, 0, 1378598912, -1677718799, 2},{0, 0, 0, 0, 0, 0, 164, 0, 0, 0, -1744830464, 2},{201392128, 0, 402653184, 2218088, 0, 0, 700448935, 675840, 0, 0, 0, 0},{0, 49169, 0, 0, 0, 0, 801112064, 1468006400, -1090518276, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 822083584, 0, 0, 0, 2656, 0},{256, 0, 20480, 0, 1275068416, 667176, 123, 0, 0, 0, -201326592, 1},{0, 0, 0, 0, 0, 255852544, 166, 0, -1073741064, 2013265920, -268432799, 1},{0, 0, 0, 0, 2016081408, 738199, 822083782, 0, 0, 0, -268435456, 1},{0, 0, 0, 0, 0, 1328512, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 696254464, 0, -1442840576, 0, 2784, 0},{262464, 0, 24576, 1879048192, 1278793809, 1322524, 692060325, 0, 0, 0, -1677721600, 2},{0, 0, 0, 0, 0, 0, 696590500, 696320, -1442839880, 1546354688, -1744827775, 2},{0, 0, 0, -1543503872, 1448151669, 738327, 796917924, 778240, -1107296256, 0, -1744830464, 2},{0, 0, 0, 0, 1761607680, 935197, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{64, 0, 0, 0, 0, 0, 197, 0, 0, 2768896, 0, 0},{0, 0, 0, 0, 0, 0, 696590336, 0, -1107296256, 0, 0, 0},{0, 0, 0, 0, 1350565888, 1353885, 0, 0, -1056964608, 0, 0, 0},{0, 0, 0, 0, 0, 0, 199, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{131072, 49168, 0, 0, 0, 0, 717225984, 0, -1358953812, 0, -1543503872, 2},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{201326592, 16777216, 8, 0, 0, 0, 0, 700416, 700, 2867200, 2704, 0},{67108864, 0, 0, 0, 0, 0, 801112064, 782336, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 2752512, -1610610048, 2},{0, 16, 0, 8398860, 0, 0, 167, 0, 764, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 196, 0, 680, 2850816, 0, 0},{0, 100663296, 16404, 1879048192, 1278269617, 1062444, 0, 0, 0, 2768896, -1543501168, 2},{0, 0, 0, 0, 0, 0, 713031680, 1460314112, -1375731032, 2850816, -1610610048, 2},{0, 0, 0, 603979776, -2025761662, 411849816, 796917958, 778240, -1073741064, 2752512, -1610610048, 2},{0, 0, 0, 603979776, -884910974, 1074094, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{131072, 0, 140, 0, 0, 0, 734003200, 0, 0, 0, -1268544400, 2},{0, 0, 0, 0, 0, 0, 170, 0, 0, 0, -1342177280, 2},{201326592, 16384, 402653184, 2218088, 0, 0, 0, 700416, -1358953796, 0, 0, 0},{201457728, 0, 0, 0, 0, 0, 801112263, 782336, -1056964608, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 720896, -1375731712, 0, 402653184, 3},{262464, 0, 24576, 1879048192, 1279842369, 929316, 717226155, 0, 0, 0, -1275068416, 2},{0, 0, 0, 0, 0, 356515840, 713388208, 720896, -1375731016, 0, -1335686048, 2},{0, 0, 0, 536870912, 1161368949, 1228179, 797266118, 778240, -1073741824, 0, 408289280, 3},{0, 0, 0, 0, -1689603072, 357714832, 190, 778240, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1228160, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{65536, 50331648, 8192, 0, 0, 0, 742391808, 716800, 0, 3260416, -872415232, 2},{0, 0, 0, 0, 0, 0, 0, 712704, 0, 0, 0, 0},{0, 48, 4, 18974816, 0, 0, 177, 0, 700, 0, 3184, 0},{131136, 0, 0, 0, 0, 0, 801112263, 0, -1056964608, 0, 0, 0},{0, 0, 0, 0, 0, 0, 191, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{268763136, 0, 0, 0, 0, 0, 734003200, 716800, 0, 0, 0, 0},{0, 0, 0, 0, 0, 415236096, 738554032, 712704, 0, 3244032, -939520928, 2},{0, 0, 0, -1409286144, 642951332, 699861, 797274302, 712704, -1073741824, 0, 0, 0},{0, 0, 0, 0, 721420288, 1354665, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{6, 16777216, 0, 2195456, 0, 371195904, 199, 0, 0, 3260416, 0, 0},{64, 0, 0, 0, 0, 0, 191, 0, -1056964608, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 16384, 0, 0, 0, 0, 0, 0, 0, -872415232, 2},{0, 0, 0, 0, 0, 398458880, 198, 0, -1073741824, 3244032, -939524096, 2},{0, 0, 0, 0, -1962934272, 1524632, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 536873984, 3},{64, 0, 0, 8421696, 0, 0, 199, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 81920, 16384, 0, 0, 0, 0, 0, -1056964608, 0, 603979776, 3},{0, 0, 0, 0, 0, 0, 200, 0, 0, 0, 677642240, 3},{0, 0, 0, 0, 0, 1460736, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 738197504, 3},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}};

//For 1st BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_A_addr;
reg [31:0]bram_ZYNQ_block_A_din;
wire [31:0]bram_ZYNQ_block_A_dout;
wire bram_ZYNQ_block_A_en;
wire [3:0]bram_ZYNQ_block_A_we;

//For 2nd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_B_addr;
reg [31:0]bram_ZYNQ_block_B_din;
wire [31:0]bram_ZYNQ_block_B_dout;
wire bram_ZYNQ_block_B_en;
wire [3:0]bram_ZYNQ_block_B_we;

//For 3rd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_C_addr;
reg [31:0]bram_ZYNQ_block_C_din;
wire [31:0]bram_ZYNQ_block_C_dout;
wire bram_ZYNQ_block_C_en;
wire [3:0]bram_ZYNQ_block_C_we;

//For 4th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_D_addr;
reg [31:0]bram_ZYNQ_block_D_din;
wire [31:0]bram_ZYNQ_block_D_dout;
wire bram_ZYNQ_block_D_en;
wire [3:0]bram_ZYNQ_block_D_we;

//For 5th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_E_addr;
reg [31:0]bram_ZYNQ_block_E_din;
wire [31:0]bram_ZYNQ_block_E_dout;
wire bram_ZYNQ_block_E_en;
wire [3:0]bram_ZYNQ_block_E_we;

//For 6th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_F_addr;
reg [31:0]bram_ZYNQ_block_F_din;
wire [31:0]bram_ZYNQ_block_F_dout;
wire bram_ZYNQ_block_F_en;
wire [3:0]bram_ZYNQ_block_F_we;

//For 7th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_G_addr;
reg [31:0]bram_ZYNQ_block_G_din;
wire [31:0]bram_ZYNQ_block_G_dout;
wire bram_ZYNQ_block_G_en;
wire [3:0]bram_ZYNQ_block_G_we;

//For 8th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_H_addr;
reg [31:0]bram_ZYNQ_block_H_din;
wire [31:0]bram_ZYNQ_block_H_dout;
wire bram_ZYNQ_block_H_en;
wire [3:0]bram_ZYNQ_block_H_we;

//Instruction BRAM
wire [31:0]bram_ZYNQ_INST_addr;
wire bram_ZYNQ_INST_en;
wire bram_ZYNQ_INST_we;

wire [31:0]bram_ZYNQ_INST_din_part_0;
wire [31:0]bram_ZYNQ_INST_din_part_1;
wire [31:0]bram_ZYNQ_INST_din_part_2;
wire [31:0]bram_ZYNQ_INST_din_part_3;
wire [31:0]bram_ZYNQ_INST_din_part_4;
wire [31:0]bram_ZYNQ_INST_din_part_5;
wire [31:0]bram_ZYNQ_INST_din_part_6;
wire [31:0]bram_ZYNQ_INST_din_part_7;
wire [31:0]bram_ZYNQ_INST_din_part_8;
wire [31:0]bram_ZYNQ_INST_din_part_9;
wire [31:0]bram_ZYNQ_INST_din_part_10;
wire [31:0]bram_ZYNQ_INST_din_part_11;

wire [31:0]bram_ZYNQ_INST_dout_part_0;
wire [31:0]bram_ZYNQ_INST_dout_part_1;
wire [31:0]bram_ZYNQ_INST_dout_part_2;
wire [31:0]bram_ZYNQ_INST_dout_part_3;
wire [31:0]bram_ZYNQ_INST_dout_part_4;
wire [31:0]bram_ZYNQ_INST_dout_part_5;
wire [31:0]bram_ZYNQ_INST_dout_part_6;
wire [31:0]bram_ZYNQ_INST_dout_part_7;
wire [31:0]bram_ZYNQ_INST_dout_part_8;
wire [31:0]bram_ZYNQ_INST_dout_part_9;
wire [31:0]bram_ZYNQ_INST_dout_part_10;
wire [31:0]bram_ZYNQ_INST_dout_part_11;

//debug signals
wire [1:0]debug_state;

reg [31:0]BRAM_dump[0:3][0:2047];
reg [31:0]fptr,fptr2;
integer count;
reg complete_bit;

//Mux signals for Address
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_dout;
reg [1:0]sel_mux_dataBRAM;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_E_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_F_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_G_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_H_dout;

//Mux signals for enable
reg mux_dataBRAM_A_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_en1 = 0; //For clearing
reg mux_dataBRAM_A_en2 = 0; //For loading A matrix
reg mux_dataBRAM_A_en3 = 0; //Currently unused
wire mux_dataBRAM_A_endout;

reg mux_dataBRAM_B_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_en1 = 0; //For clearing
reg mux_dataBRAM_B_en2 = 0; //For loading A matrix
reg mux_dataBRAM_B_en3 = 0; //Currently unused
wire mux_dataBRAM_B_endout;

reg mux_dataBRAM_C_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_en1 = 0; //For clearing
reg mux_dataBRAM_C_en2 = 0; //For loading A matrix
reg mux_dataBRAM_C_en3 = 0; //Currently unused
wire mux_dataBRAM_C_endout;

reg mux_dataBRAM_D_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_en1 = 0; //For clearing
reg mux_dataBRAM_D_en2 = 0; //For loading A matrix
reg mux_dataBRAM_D_en3 = 0; //Currently unused
wire mux_dataBRAM_D_endout;

reg mux_dataBRAM_E_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_E_en1 = 0; //For clearing
reg mux_dataBRAM_E_en2 = 0; //For loading A matrix
reg mux_dataBRAM_E_en3 = 0; //Currently unused
wire mux_dataBRAM_E_endout;

reg mux_dataBRAM_F_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_F_en1 = 0; //For clearing
reg mux_dataBRAM_F_en2 = 0; //For loading A matrix
reg mux_dataBRAM_F_en3 = 0; //Currently unused
wire mux_dataBRAM_F_endout;

reg mux_dataBRAM_G_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_G_en1 = 0; //For clearing
reg mux_dataBRAM_G_en2 = 0; //For loading A matrix
reg mux_dataBRAM_G_en3 = 0; //Currently unused
wire mux_dataBRAM_G_endout;

reg mux_dataBRAM_H_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_H_en1 = 0; //For clearing
reg mux_dataBRAM_H_en2 = 0; //For loading A matrix
reg mux_dataBRAM_H_en3 = 0; //Currently unused
wire mux_dataBRAM_H_endout;

//Mux signals for write enable
reg mux_dataBRAM_A_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_we1 = 0; //For clearing
reg mux_dataBRAM_A_we2 = 0; //For loading A matrix
reg mux_dataBRAM_A_we3 = 0; //Currently unused
wire mux_dataBRAM_A_wedout;

reg mux_dataBRAM_B_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_we1 = 0; //For clearing
reg mux_dataBRAM_B_we2 = 0; //For loading A matrix
reg mux_dataBRAM_B_we3 = 0; //Currently unused
wire mux_dataBRAM_B_wedout;

reg mux_dataBRAM_C_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_we1 = 0; //For clearing
reg mux_dataBRAM_C_we2 = 0; //For loading A matrix
reg mux_dataBRAM_C_we3 = 0; //Currently unused
wire mux_dataBRAM_C_wedout;

reg mux_dataBRAM_D_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_we1 = 0; //For clearing
reg mux_dataBRAM_D_we2 = 0; //For loading A matrix
reg mux_dataBRAM_D_we3 = 0; //Currently unused
wire mux_dataBRAM_D_wedout;

reg mux_dataBRAM_E_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_E_we1 = 0; //For clearing
reg mux_dataBRAM_E_we2 = 0; //For loading A matrix
reg mux_dataBRAM_E_we3 = 0; //Currently unused
wire mux_dataBRAM_E_wedout;

reg mux_dataBRAM_F_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_F_we1 = 0; //For clearing
reg mux_dataBRAM_F_we2 = 0; //For loading A matrix
reg mux_dataBRAM_F_we3 = 0; //Currently unused
wire mux_dataBRAM_F_wedout;

reg mux_dataBRAM_G_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_G_we1 = 0; //For clearing
reg mux_dataBRAM_G_we2 = 0; //For loading A matrix
reg mux_dataBRAM_G_we3 = 0; //Currently unused
wire mux_dataBRAM_G_wedout;

reg mux_dataBRAM_H_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_H_we1 = 0; //For clearing
reg mux_dataBRAM_H_we2 = 0; //For loading A matrix
reg mux_dataBRAM_H_we3 = 0; //Currently unused
wire mux_dataBRAM_H_wedout;

//Mux signals for din
reg [31:0]mux_dataBRAM_A_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_A_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_A_din_out;
reg sel_mux_dataBRAM_din;

reg [31:0]mux_dataBRAM_B_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_B_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_B_din_out;

reg [31:0]mux_dataBRAM_C_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_C_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_C_din_out;

reg [31:0]mux_dataBRAM_D_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_D_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_D_din_out;

reg [31:0]mux_dataBRAM_E_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_E_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_E_din_out;

reg [31:0]mux_dataBRAM_F_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_F_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_F_din_out;

reg [31:0]mux_dataBRAM_G_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_G_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_G_din_out;

reg [31:0]mux_dataBRAM_H_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_H_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_H_din_out;

//Instruction BRAM muxes
reg [31:0]instBRAM_part0_din;
reg [31:0]instBRAM_part1_din;
reg [31:0]instBRAM_part2_din;
reg [31:0]instBRAM_part3_din;
reg [31:0]instBRAM_part4_din;
reg [31:0]instBRAM_part5_din;
reg [31:0]instBRAM_part6_din;
reg [31:0]instBRAM_part7_din;
reg [31:0]instBRAM_part8_din;
reg [31:0]instBRAM_part9_din;
reg [31:0]instBRAM_part10_din;
reg [31:0]instBRAM_part11_din;

reg instBRAM_en = 0;
reg instBRAM_we = 0;
reg [ADDR_WIDTH-1:0]instBRAM_addr;


//Memory dump start and complete signals
reg start_mem_dump;
reg mem_dump_complete;
reg start_dataBRAM_erase;
reg dataBRAM_erase_complete;
reg start_A_load;
reg A_load_complete;
reg start_instBRAM_erase;
reg instBRAM_erase_complete;
reg start_inst_load;
reg inst_load_complete;
reg start_full_run;
reg complete_full_run;
reg start0; //For full run
reg complete_sig;

LUDH_TEST_WRAPPER #(ADDR_WIDTH,ADDR_WIDTH_DATA_BRAM,CTRL_WIDTH,AU_SEL_WIDTH,BRAM_SEL_WIDTH) uut1 (
CLK_100,

locked,
RST_IN,
start_sig,
completed,

//First BRAM
bram_ZYNQ_block_A_addr, 
bram_ZYNQ_block_A_din, 
bram_ZYNQ_block_A_dout, 
bram_ZYNQ_block_A_en,
bram_ZYNQ_block_A_we, 

//Second BRAM
bram_ZYNQ_block_B_addr, 
bram_ZYNQ_block_B_din, 
bram_ZYNQ_block_B_dout, 
bram_ZYNQ_block_B_en,
bram_ZYNQ_block_B_we, 

//Third BRAM
bram_ZYNQ_block_C_addr, 
bram_ZYNQ_block_C_din, 
bram_ZYNQ_block_C_dout, 
bram_ZYNQ_block_C_en,
bram_ZYNQ_block_C_we, 

//Fourth BRAM
bram_ZYNQ_block_D_addr, 
bram_ZYNQ_block_D_din, 
bram_ZYNQ_block_D_dout, 
bram_ZYNQ_block_D_en,
bram_ZYNQ_block_D_we, 

//Fifth BRAM
bram_ZYNQ_block_E_addr, 
bram_ZYNQ_block_E_din, 
bram_ZYNQ_block_E_dout, 
bram_ZYNQ_block_E_en,
bram_ZYNQ_block_E_we, 

//Sixth BRAM
bram_ZYNQ_block_F_addr, 
bram_ZYNQ_block_F_din, 
bram_ZYNQ_block_F_dout, 
bram_ZYNQ_block_F_en,
bram_ZYNQ_block_F_we, 

//Seventh BRAM
bram_ZYNQ_block_G_addr, 
bram_ZYNQ_block_G_din, 
bram_ZYNQ_block_G_dout, 
bram_ZYNQ_block_G_en,
bram_ZYNQ_block_G_we, 

//Eighth BRAM
bram_ZYNQ_block_H_addr, 
bram_ZYNQ_block_H_din, 
bram_ZYNQ_block_H_dout, 
bram_ZYNQ_block_H_en,
bram_ZYNQ_block_H_we, 

//Instruction BRAM
bram_ZYNQ_INST_addr,
bram_ZYNQ_INST_en,
bram_ZYNQ_INST_we,
        
bram_ZYNQ_INST_din_part_0,
bram_ZYNQ_INST_din_part_1,
bram_ZYNQ_INST_din_part_2,
bram_ZYNQ_INST_din_part_3,
bram_ZYNQ_INST_din_part_4,
bram_ZYNQ_INST_din_part_5,
bram_ZYNQ_INST_din_part_6,
bram_ZYNQ_INST_din_part_7,
bram_ZYNQ_INST_din_part_8,
bram_ZYNQ_INST_din_part_9,
bram_ZYNQ_INST_din_part_10,
bram_ZYNQ_INST_din_part_11,
        
bram_ZYNQ_INST_dout_part_0,
bram_ZYNQ_INST_dout_part_1,
bram_ZYNQ_INST_dout_part_2,
bram_ZYNQ_INST_dout_part_3,
bram_ZYNQ_INST_dout_part_4,
bram_ZYNQ_INST_dout_part_5,
bram_ZYNQ_INST_dout_part_6,
bram_ZYNQ_INST_dout_part_7,
bram_ZYNQ_INST_dout_part_8,
bram_ZYNQ_INST_dout_part_9,
bram_ZYNQ_INST_dout_part_10,
bram_ZYNQ_INST_dout_part_11,
        
//debug signals
debug_state
);

initial begin
CLK_100 = 1'b1;
forever #(t_100/2) CLK_100 = ~CLK_100;
end

//Initiallizing the mux to be used for DATA BRAMS address multiplexing
//For address
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut2(mux_dataBRAM_A_dout,mux_dataBRAM_A_0,mux_dataBRAM_A_1,mux_dataBRAM_A_2,mux_dataBRAM_A_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut3(mux_dataBRAM_B_dout,mux_dataBRAM_B_0,mux_dataBRAM_B_1,mux_dataBRAM_B_2,mux_dataBRAM_B_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut4(mux_dataBRAM_C_dout,mux_dataBRAM_C_0,mux_dataBRAM_C_1,mux_dataBRAM_C_2,mux_dataBRAM_C_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut5(mux_dataBRAM_D_dout,mux_dataBRAM_D_0,mux_dataBRAM_D_1,mux_dataBRAM_D_2,mux_dataBRAM_D_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut18(mux_dataBRAM_E_dout,mux_dataBRAM_E_0,mux_dataBRAM_E_1,mux_dataBRAM_E_2,mux_dataBRAM_E_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut19(mux_dataBRAM_F_dout,mux_dataBRAM_F_0,mux_dataBRAM_F_1,mux_dataBRAM_F_2,mux_dataBRAM_F_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut20(mux_dataBRAM_G_dout,mux_dataBRAM_G_0,mux_dataBRAM_G_1,mux_dataBRAM_G_2,mux_dataBRAM_G_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut21(mux_dataBRAM_H_dout,mux_dataBRAM_H_0,mux_dataBRAM_H_1,mux_dataBRAM_H_2,mux_dataBRAM_H_3,sel_mux_dataBRAM);

//For enable
mux_4x1 #(1) uut6(mux_dataBRAM_A_endout,mux_dataBRAM_A_en0,mux_dataBRAM_A_en1,mux_dataBRAM_A_en2,mux_dataBRAM_A_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut7(mux_dataBRAM_B_endout,mux_dataBRAM_B_en0,mux_dataBRAM_B_en1,mux_dataBRAM_B_en2,mux_dataBRAM_B_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut8(mux_dataBRAM_C_endout,mux_dataBRAM_C_en0,mux_dataBRAM_C_en1,mux_dataBRAM_C_en2,mux_dataBRAM_C_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut9(mux_dataBRAM_D_endout,mux_dataBRAM_D_en0,mux_dataBRAM_D_en1,mux_dataBRAM_D_en2,mux_dataBRAM_D_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut22(mux_dataBRAM_E_endout,mux_dataBRAM_E_en0,mux_dataBRAM_E_en1,mux_dataBRAM_E_en2,mux_dataBRAM_E_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut23(mux_dataBRAM_F_endout,mux_dataBRAM_F_en0,mux_dataBRAM_F_en1,mux_dataBRAM_F_en2,mux_dataBRAM_F_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut24(mux_dataBRAM_G_endout,mux_dataBRAM_G_en0,mux_dataBRAM_G_en1,mux_dataBRAM_G_en2,mux_dataBRAM_G_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut25(mux_dataBRAM_H_endout,mux_dataBRAM_H_en0,mux_dataBRAM_H_en1,mux_dataBRAM_H_en2,mux_dataBRAM_H_en3,sel_mux_dataBRAM);

//For Write enable
mux_4x1 #(1) uut10(mux_dataBRAM_A_wedout,mux_dataBRAM_A_we0,mux_dataBRAM_A_we1,mux_dataBRAM_A_we2,mux_dataBRAM_A_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut11(mux_dataBRAM_B_wedout,mux_dataBRAM_B_we0,mux_dataBRAM_B_we1,mux_dataBRAM_B_we2,mux_dataBRAM_B_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut12(mux_dataBRAM_C_wedout,mux_dataBRAM_C_we0,mux_dataBRAM_C_we1,mux_dataBRAM_C_we2,mux_dataBRAM_C_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut13(mux_dataBRAM_D_wedout,mux_dataBRAM_D_we0,mux_dataBRAM_D_we1,mux_dataBRAM_D_we2,mux_dataBRAM_D_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut26(mux_dataBRAM_E_wedout,mux_dataBRAM_E_we0,mux_dataBRAM_E_we1,mux_dataBRAM_E_we2,mux_dataBRAM_E_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut27(mux_dataBRAM_F_wedout,mux_dataBRAM_F_we0,mux_dataBRAM_F_we1,mux_dataBRAM_F_we2,mux_dataBRAM_F_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut28(mux_dataBRAM_G_wedout,mux_dataBRAM_G_we0,mux_dataBRAM_G_we1,mux_dataBRAM_G_we2,mux_dataBRAM_G_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut29(mux_dataBRAM_H_wedout,mux_dataBRAM_H_we0,mux_dataBRAM_H_we1,mux_dataBRAM_H_we2,mux_dataBRAM_H_we3,sel_mux_dataBRAM);

//For din
mux_2x1 #(32) uut14(mux_dataBRAM_A_din_out,mux_dataBRAM_A_din0,mux_dataBRAM_A_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut15(mux_dataBRAM_B_din_out,mux_dataBRAM_B_din0,mux_dataBRAM_B_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut16(mux_dataBRAM_C_din_out,mux_dataBRAM_C_din0,mux_dataBRAM_C_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut17(mux_dataBRAM_D_din_out,mux_dataBRAM_D_din0,mux_dataBRAM_D_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut30(mux_dataBRAM_E_din_out,mux_dataBRAM_E_din0,mux_dataBRAM_E_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut31(mux_dataBRAM_F_din_out,mux_dataBRAM_F_din0,mux_dataBRAM_F_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut32(mux_dataBRAM_G_din_out,mux_dataBRAM_G_din0,mux_dataBRAM_G_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut33(mux_dataBRAM_H_din_out,mux_dataBRAM_H_din0,mux_dataBRAM_H_din1,sel_mux_dataBRAM_din);


initial begin
start_mem_dump <= 0;
mem_dump_complete <= 0;
start_dataBRAM_erase <= 0;
dataBRAM_erase_complete <= 0;
start_A_load <= 0;
A_load_complete <= 0;
start_instBRAM_erase <= 0;
instBRAM_erase_complete <= 0;
start_inst_load <= 0;
inst_load_complete <= 0;
complete_full_run <= 0;
sel_mux_dataBRAM <= 2'b00;
sel_mux_dataBRAM_din <= 1'b0;

count <= -1;
complete_bit <= 1'b0;
locked <= 1'b0;

#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
RST_IN <= 1'b1;

//Resetting the contents of data BRAMS and Inst BRAM
#(t_100*50)
sel_mux_dataBRAM <= 2'b01;
sel_mux_dataBRAM_din <= 1'b0;
start_dataBRAM_erase <= 1'b1;

@(posedge dataBRAM_erase_complete)
#(t_100*50)
start_dataBRAM_erase <= 0;

#(t_100*50)
start_instBRAM_erase <= 1'b1;

@(posedge instBRAM_erase_complete)
#(t_100*50)
start_instBRAM_erase <= 0;

//Loading the A matrix
#(t_100*50)
sel_mux_dataBRAM <= 2'b10;
sel_mux_dataBRAM_din <= 1'b1;
start_A_load <= 1'b1;

@(posedge A_load_complete)
#(t_100*50)
start_A_load <= 0;

//RST = 0
#(t_100*50)
RST_IN <= 1'b0;

//Locked = 1
#(t_100*50)
locked <= 1'b1;

//Loading the instruction matrix and starting LU Decomposition
#(t_100*50)
start_full_run = 1'b1;

@(posedge complete_sig)
complete_bit <= 1'b1;
#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
sel_mux_dataBRAM <= 2'b00;
start_mem_dump <= 1;

@(posedge mem_dump_complete)
#(t_100*50)
start_mem_dump <= 0;
$stop;

end

assign start_sig = start0;
assign complete_sig = complete_full_run;

//Address signals(data BRAM)
assign bram_ZYNQ_block_A_addr = mux_dataBRAM_A_dout;
assign bram_ZYNQ_block_B_addr = mux_dataBRAM_B_dout;
assign bram_ZYNQ_block_C_addr = mux_dataBRAM_C_dout;
assign bram_ZYNQ_block_D_addr = mux_dataBRAM_D_dout;
assign bram_ZYNQ_block_E_addr = mux_dataBRAM_E_dout;
assign bram_ZYNQ_block_F_addr = mux_dataBRAM_F_dout;
assign bram_ZYNQ_block_G_addr = mux_dataBRAM_G_dout;
assign bram_ZYNQ_block_H_addr = mux_dataBRAM_H_dout;

//Enable signals(data BRAM)
assign bram_ZYNQ_block_A_en = mux_dataBRAM_A_endout;
assign bram_ZYNQ_block_B_en = mux_dataBRAM_B_endout;
assign bram_ZYNQ_block_C_en = mux_dataBRAM_C_endout;
assign bram_ZYNQ_block_D_en = mux_dataBRAM_D_endout;
assign bram_ZYNQ_block_E_en = mux_dataBRAM_E_endout;
assign bram_ZYNQ_block_F_en = mux_dataBRAM_F_endout;
assign bram_ZYNQ_block_G_en = mux_dataBRAM_G_endout;
assign bram_ZYNQ_block_H_en = mux_dataBRAM_H_endout;

//Write enable signals(data BRAM)
assign bram_ZYNQ_block_A_we = mux_dataBRAM_A_wedout;
assign bram_ZYNQ_block_B_we = mux_dataBRAM_B_wedout;
assign bram_ZYNQ_block_C_we = mux_dataBRAM_C_wedout;
assign bram_ZYNQ_block_D_we = mux_dataBRAM_D_wedout;
assign bram_ZYNQ_block_E_we = mux_dataBRAM_E_wedout;
assign bram_ZYNQ_block_F_we = mux_dataBRAM_F_wedout;
assign bram_ZYNQ_block_G_we = mux_dataBRAM_G_wedout;
assign bram_ZYNQ_block_H_we = mux_dataBRAM_H_wedout;

//din signals(data BRAM)
assign bram_ZYNQ_block_A_din = mux_dataBRAM_A_din_out;
assign bram_ZYNQ_block_B_din = mux_dataBRAM_B_din_out;
assign bram_ZYNQ_block_C_din = mux_dataBRAM_C_din_out;
assign bram_ZYNQ_block_D_din = mux_dataBRAM_D_din_out;
assign bram_ZYNQ_block_E_din = mux_dataBRAM_E_din_out;
assign bram_ZYNQ_block_F_din = mux_dataBRAM_F_din_out;
assign bram_ZYNQ_block_G_din = mux_dataBRAM_G_din_out;
assign bram_ZYNQ_block_H_din = mux_dataBRAM_H_din_out;

//Address signal(inst BRAM)
assign bram_ZYNQ_INST_addr = instBRAM_addr;

//Enable signal(inst BRAM)
assign bram_ZYNQ_INST_en = instBRAM_en;

//Write enable signal(inst BRAM)
assign bram_ZYNQ_INST_we = instBRAM_we;

//din signal(inst BRAM)
assign bram_ZYNQ_INST_din_part_0 = instBRAM_part0_din;
assign bram_ZYNQ_INST_din_part_1 = instBRAM_part1_din;
assign bram_ZYNQ_INST_din_part_2 = instBRAM_part2_din;
assign bram_ZYNQ_INST_din_part_3 = instBRAM_part3_din;
assign bram_ZYNQ_INST_din_part_4 = instBRAM_part4_din;
assign bram_ZYNQ_INST_din_part_5 = instBRAM_part5_din;
assign bram_ZYNQ_INST_din_part_6 = instBRAM_part6_din;
assign bram_ZYNQ_INST_din_part_7 = instBRAM_part7_din;
assign bram_ZYNQ_INST_din_part_8 = instBRAM_part8_din;
assign bram_ZYNQ_INST_din_part_9 = instBRAM_part9_din;
assign bram_ZYNQ_INST_din_part_10 = instBRAM_part10_din;
assign bram_ZYNQ_INST_din_part_11 = instBRAM_part11_din;


//Always block for full run
always@(posedge CLK_100) begin
if(CLK_100  == 1 && start_full_run == 1 && complete_full_run != 1) begin
//Start loading complete instructions
start_inst_load <= 1'b1;
@(posedge inst_load_complete)
#(t_100*50)
start_inst_load <= 0;

//Start the LU Decomposition
#(t_100*50)
start0 <= 1'b1;
complete_full_run <= 1'b0;

//Waiting for completion
@(posedge completed)
complete_full_run <= 1'b1;

end
else if(CLK_100 == 1 && start_full_run == 0) begin
start0 <= 0;
complete_full_run <= 0;
end
end

//Always block to dump bram contents
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_mem_dump == 1 && mem_dump_complete != 1)begin 

    if(count == -1) begin
        fptr = $fopen("BRAM_dump.txt","w");
        $fdisplay(fptr,"float bram_dump[%d][%d];",BRAM_LIMIT_IND_DEBUG,DATA_BRAM_SIZE);
        mux_dataBRAM_A_en0 = 1'b1; mux_dataBRAM_B_en0 = 1'b1; mux_dataBRAM_C_en0 = 1'b1; mux_dataBRAM_D_en0 = 1'b1; mux_dataBRAM_E_en0 = 1'b1; mux_dataBRAM_F_en0 = 1'b1; mux_dataBRAM_G_en0 = 1'b1; mux_dataBRAM_H_en0 = 1'b1;
        mux_dataBRAM_A_we0 = 1'b0; mux_dataBRAM_B_we0 = 1'b0; mux_dataBRAM_C_we0 = 1'b0; mux_dataBRAM_D_we0 = 1'b0; mux_dataBRAM_E_we0 = 1'b0; mux_dataBRAM_F_we0 = 1'b0; mux_dataBRAM_G_we0 = 1'b0; mux_dataBRAM_H_we0 = 1'b0;
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];
    end
    else if(count == 0) begin
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Addres
    end
    else if(count <= DATA_BRAM_SIZE && count >= 1)begin
        $fdisplay(fptr,"bram_dump[0][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_A_dout)); //count-1 because BRAM has single cycle latency
        $fdisplay(fptr,"bram_dump[1][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_B_dout));
        $fdisplay(fptr,"bram_dump[2][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_C_dout));
        $fdisplay(fptr,"bram_dump[3][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_D_dout));
        $fdisplay(fptr,"bram_dump[4][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_E_dout));
        $fdisplay(fptr,"bram_dump[5][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_F_dout));
        $fdisplay(fptr,"bram_dump[6][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_G_dout));
        $fdisplay(fptr,"bram_dump[7][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_H_dout));
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Address
    end
    else if (count == DATA_BRAM_SIZE+1) begin
        $fclose(fptr);
        count = -1;
        mem_dump_complete = 1;    
        mux_dataBRAM_A_en0 = 1'b0; mux_dataBRAM_B_en0 = 1'b0; mux_dataBRAM_C_en0 = 1'b0; mux_dataBRAM_D_en0 = 1'b0; mux_dataBRAM_E_en0 = 1'b0; mux_dataBRAM_F_en0 = 1'b0; mux_dataBRAM_G_en0 = 1'b0; mux_dataBRAM_H_en0 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_mem_dump == 0)
    mem_dump_complete = 0;
end


//Always block to erase data BRAM contents
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_dataBRAM_erase == 1 && dataBRAM_erase_complete != 1)begin 

    if(count <= DATA_BRAM_SIZE-2 && count >= -1)begin
        if(count == -1) begin
            mux_dataBRAM_A_en1 = 1'b1; mux_dataBRAM_B_en1 = 1'b1; mux_dataBRAM_C_en1 = 1'b1; mux_dataBRAM_D_en1 = 1'b1; mux_dataBRAM_E_en1 = 1'b1; mux_dataBRAM_F_en1 = 1'b1; mux_dataBRAM_G_en1 = 1'b1; mux_dataBRAM_H_en1 = 1'b1;
            mux_dataBRAM_A_we1 = 1'b1; mux_dataBRAM_B_we1 = 1'b1; mux_dataBRAM_C_we1 = 1'b1; mux_dataBRAM_D_we1 = 1'b1; mux_dataBRAM_E_we1 = 1'b1; mux_dataBRAM_F_we1 = 1'b1; mux_dataBRAM_G_we1 = 1'b1; mux_dataBRAM_H_we1 = 1'b1;
            mux_dataBRAM_A_din0 = 0; mux_dataBRAM_B_din0 = 0; mux_dataBRAM_C_din0 = 0; mux_dataBRAM_D_din0 = 0; mux_dataBRAM_E_din0 = 0; mux_dataBRAM_F_din0 = 0; mux_dataBRAM_G_din0 = 0; mux_dataBRAM_H_din0 = 0; //Reset value
        end
        count = count + 1;
        mux_dataBRAM_A_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_E_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_F_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_G_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_H_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; //Address
    end
    else if (count == DATA_BRAM_SIZE-1) begin
        count = -1;
        dataBRAM_erase_complete = 1;   
        mux_dataBRAM_A_en1 = 1'b0; mux_dataBRAM_B_en1 = 1'b0; mux_dataBRAM_C_en1 = 1'b0; mux_dataBRAM_D_en1 = 1'b0; mux_dataBRAM_E_en1 = 1'b0; mux_dataBRAM_F_en1 = 1'b0; mux_dataBRAM_G_en1 = 1'b0; mux_dataBRAM_H_en1 = 1'b0;
        mux_dataBRAM_A_we1 = 1'b0; mux_dataBRAM_B_we1 = 1'b0; mux_dataBRAM_C_we1 = 1'b0; mux_dataBRAM_D_we1 = 1'b0; mux_dataBRAM_E_we1 = 1'b0; mux_dataBRAM_F_we1 = 1'b0; mux_dataBRAM_G_we1 = 1'b0; mux_dataBRAM_H_we1 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_dataBRAM_erase == 0)
    dataBRAM_erase_complete = 0;
end

//Always block to load the A matrix in data bram
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_A_load == 1 && A_load_complete != 1)begin 

    if(count <= A_size-2 && count >= -1)begin
        if(count == -1) //Initialization of en signals
            mux_dataBRAM_A_en2 = 1'b1; mux_dataBRAM_B_en2 = 1'b1; mux_dataBRAM_C_en2 = 1'b1; mux_dataBRAM_D_en2 = 1'b1; mux_dataBRAM_E_en2 = 1'b1; mux_dataBRAM_F_en2 = 1'b1; mux_dataBRAM_G_en2 = 1'b1; mux_dataBRAM_H_en2 = 1'b1;
            
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0; mux_dataBRAM_E_we2 = 1'b0; mux_dataBRAM_F_we2 = 1'b0; mux_dataBRAM_G_we2 = 1'b0; mux_dataBRAM_H_we2 = 1'b0;//Initially assigning all the write enables to 0
        count = count + 1;
        if(A_BRAMInd[count] == 0) begin//making one of the write enables 1
            mux_dataBRAM_A_we2 = 1'b1; mux_dataBRAM_A_2 = A_BRAMAddr[count]; mux_dataBRAM_A_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 1) begin
            mux_dataBRAM_B_we2 = 1'b1; mux_dataBRAM_B_2 = A_BRAMAddr[count]; mux_dataBRAM_B_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 2) begin
            mux_dataBRAM_C_we2 = 1'b1; mux_dataBRAM_C_2 = A_BRAMAddr[count]; mux_dataBRAM_C_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 3) begin
            mux_dataBRAM_D_we2 = 1'b1; mux_dataBRAM_D_2 = A_BRAMAddr[count]; mux_dataBRAM_D_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 4) begin
            mux_dataBRAM_E_we2 = 1'b1; mux_dataBRAM_E_2 = A_BRAMAddr[count]; mux_dataBRAM_E_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 5) begin
            mux_dataBRAM_F_we2 = 1'b1; mux_dataBRAM_F_2 = A_BRAMAddr[count]; mux_dataBRAM_F_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 6) begin
            mux_dataBRAM_G_we2 = 1'b1; mux_dataBRAM_G_2 = A_BRAMAddr[count]; mux_dataBRAM_G_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 7) begin
            mux_dataBRAM_H_we2 = 1'b1; mux_dataBRAM_H_2 = A_BRAMAddr[count]; mux_dataBRAM_H_din1 = A[count];
        end
    end
    else if (count == A_size-1) begin
        count = -1;
        A_load_complete = 1;   
        mux_dataBRAM_A_en2 = 1'b0; mux_dataBRAM_B_en2 = 1'b0; mux_dataBRAM_C_en2 = 1'b0; mux_dataBRAM_D_en2 = 1'b0; mux_dataBRAM_E_en2 = 1'b0; mux_dataBRAM_F_en2 = 1'b0; mux_dataBRAM_G_en2 = 1'b0; mux_dataBRAM_H_en2 = 1'b0;
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0; mux_dataBRAM_E_we2 = 1'b0; mux_dataBRAM_F_we2 = 1'b0; mux_dataBRAM_G_we2 = 1'b0; mux_dataBRAM_H_we2 = 1'b0;
    end
end
else if(CLK_100 == 1 && start_A_load == 0)
    A_load_complete = 0;
end

//Always block to erase inst BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_instBRAM_erase == 1 && instBRAM_erase_complete != 1)begin 

    if(count <= INST_BRAM_SIZE-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
            instBRAM_part0_din = 0; instBRAM_part1_din = 0; instBRAM_part2_din = 0; instBRAM_part3_din = 0; instBRAM_part4_din = 0; instBRAM_part5_din = 0;
            instBRAM_part6_din = 0; instBRAM_part7_din = 0; instBRAM_part8_din = 0; instBRAM_part9_din = 0; instBRAM_part10_din = 0; instBRAM_part11_din = 0;
        end
        count = count + 1;
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == INST_BRAM_SIZE-1) begin
        count = -1;
        instBRAM_erase_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_instBRAM_erase == 0)
    instBRAM_erase_complete = 0;
end

//Always block to load instruction to instruction BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_inst_load == 1 && inst_load_complete != 1)begin 

    if(count <= total_instructions-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
        end
        count = count + 1;
        instBRAM_part0_din = Inst[count][0]; instBRAM_part1_din = Inst[count][1]; instBRAM_part2_din = Inst[count][2]; instBRAM_part3_din = Inst[count][3]; 
        instBRAM_part4_din = Inst[count][4]; instBRAM_part5_din = Inst[count][5]; instBRAM_part6_din = Inst[count][6]; instBRAM_part7_din = Inst[count][7]; 
        instBRAM_part8_din = Inst[count][8]; instBRAM_part9_din = Inst[count][9]; instBRAM_part10_din = Inst[count][10]; instBRAM_part11_din = Inst[count][11];
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == total_instructions-1) begin
        count = -1;
        inst_load_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_inst_load == 0)
    inst_load_complete = 0;
end

function real float_conv(input [31:0]b_num);
reg sign;
reg [7:0]weighted_expt;
integer actual_expt;
reg [1:23] mantissa;
reg [7:0] i;
real temp_result,temp_decimal;

begin
sign = b_num >> 31;
weighted_expt = (b_num & 32'h7f800000)>> 23;
mantissa = b_num & 32'h007fffff;

if(weighted_expt == 0)begin
	temp_result = 1.0;
	for(i=0;i<126;i=i+1)
		temp_result = temp_result/2;

	temp_decimal = 0;
	for(i=1;i<=23;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(1.0/(1<<i));
		
	temp_result = temp_result*temp_decimal;
	if(sign==1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
	end
else if(weighted_expt>0 && weighted_expt <255) begin
	actual_expt = weighted_expt-127;
	if(actual_expt<0)begin
		temp_result = 1.0;
		actual_expt = -actual_expt;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result/2;
		end
	else begin
		temp_result = 1.0;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result*2;
	end

	temp_decimal = 0;
	for(i=1;i<=23;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(1.0/(1<<i));

	temp_decimal = temp_decimal + 1;
	temp_result = temp_result*temp_decimal;
	if(sign == 1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
end
else if(weighted_expt == 255)begin
/*if(mantissa == 0 and sign == 0)
float_conv = "inf";
else if(mantissa == 0 and sign == 1)
float_conv = "-inf";
else
float_conv = "nan";*/
end

end
endfunction

endmodule

module mux_4x1 #(parameter integer data_width = 11)(dout,din0,din1,din2,din3,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input [data_width-1:0]din2;
input [data_width-1:0]din3;
input [1:0]sel;

always@(din0,din1,din2,din3,sel) begin
case(sel)
2'b00: dout <= din0;
2'b01: dout <= din1;
2'b10: dout <= din2;
2'b11: dout <= din3;
endcase
end
endmodule

module mux_2x1 #(parameter integer data_width = 32)(dout,din0,din1,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input sel;

always@(din0,din1,sel) begin
case(sel)
1'b0: dout <= din0;
1'b1: dout <= din1;
endcase
end
endmodule













