`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.12.2019 07:59:36
// Design Name: 
// Module Name: simTester_verilog
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simTester_verilog();
reg CLK_100, CLK_200, locked, RST_IN,start_sig;
wire  completed;
localparam time t_100 = 40;
localparam time t_200 = 20;

localparam integer ADDR_WIDTH = 12;
localparam integer ADDR_WIDTH_DATA_BRAM = 11;
localparam integer CTRL_WIDTH = 373;
localparam integer AU_SEL_WIDTH = 5;
localparam integer BRAM_SEL_WIDTH = 5;

localparam integer BRAM_LIMIT_IND_DEBUG = 4; //It indicates that BRAM contents from location 0 to BRAM_LIMIT_IND_DEBUG will be dumped for all 4 BRAMS for every cycle

//Constant array to load the A matrix
localparam integer A_size = 5852;
localparam integer A[0:5851] = '{1044000396, -1578745596, -1103483252, -1646356858, 1044000396, -1416839988, -1103483252, 1044044739, -1171441730, -1103483252, -1171438918, 1044044750, -1413100403, -1103483252, 1044000396, -1399080270, -1103483252, -1449639013, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1324625067, -1103483252, -1103483252, -1382850568, 1044000396, -1416839988, -1103483252, 1044000933, -1224316244, -1416839988, -1175620078, 1044035198, -1198934101, -1103483252, 1044000680, -1232190757, -1103483252, -1303525842, 1044000396, -1416839988, -1103483252, 1065353216, 1044000680, -1232187903, -1103483252, -1303521536, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1416839988, -1103483252, 1044001095, -1221665839, -1103483252, -1103483252, -1172416790, 1044058626, -1182122023, -1103483252, 1044133849, -1157475477, -1324783727, -1157593266, 1044132009, -1416839914, -1103483252, 1044000396, -1866686131, -1103483252, -1921795428, 1044000396, -1103483252, -1416839988, 1044053186, -1169279348, -1103483252, -1168046700, 1044058024, -1263185281, -1103483252, 1044043696, -1171708920, -1103483252, -1171149725, 1044045901, -1103483252, -1263953053, 1044000396, -1103483252, -1416839988, 1044000397, -1295114178, -1103483252, -1366877434, 1044000396, -1103483252, -1416839988, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, 1044049265, -1170288757, -1263616959, -1103483252, -1103483252, -1170235283, 1044049452, -1416827917, 1044000396, -1653844636, -1103483252, -1597157163, 1044000396, -1416839988, -1103483252, 1044001666, -1214327595, -1103483252, -1173144354, 1044038100, -1271165407, -1103483252, 1044000396, 0, -1103483252, 0, 1082231448, -1065913784, -1103483252, 1065353216, -1103483252, 1044000396, -1416839988, 1044000396, -1103483252, -1103483252, 1052389004, -1103483252, -1416839988, -1103483252, 1044000396, -1774871817, -1416839988, -1717318962, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -2147467728, -1103483252, -1103483252, -2147483616, 1044000396, -1416839988, -1103483252, 1044017251, -1182552145, -1416839988, -1183913376, 1044015686, -1416839988, -1103483252, 1065353216, -1103483251, 1044042947, -1171900841, -1416839198, -1172369804, 1044041114, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044083025, -1163828580, -1350897415, -1103483252, -1163860672, 1044082774, -1065913784, -1103483252, 1082231448, -1307130875, -1416839988, -1362934801, 1044000396, -1103483252, -1103483252, 1044050074, -1170075973, -1236687943, -1170121374, 1044050099, -1103483252, -1103483252, 1044000396, -2147483593, -1416839988, 0, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044032013, -1174994422, -1416839988, -1103483252, -1183875328, 1044015723, -1186107103, -1103483252, 1044044743, -1175208367, -1416839988, -1184998193, 1044014627, -1103483252, -1103483252, -1103483252, -1187663181, 959820467, 1052389004, -1103483252, -1103483252, -1310599885, 836883763, -1186124833, 961358815, 1052389004, 550205209, -1597278439, 971952289, -1175531359, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103489106, -1195946757, -1103483252, -1416839988, -1416839988, -1416839988, 1063831305, -1103482052, 932568763, -1103483252, -1416839988, -1103478592, 949068995, -1182485878, 946851788, 1065353216, -1103483252, -1416839988, -1103483252, -1065913784, 1091192010, -1103483252, -1416839988, -1416839988, -1416839988, -1103483206, 892907363, -1065913784, 823212534, -1103483208, -1239626935, 1065353216, 935366344, -1212117304, -1297403033, 850080615, -1103483252, -1103483252, 1052389004, -1103483252, -1103483252, -2147473575, 10073, -1236498597, 910985051, -1241218894, 906264754, -2147483614, 34, 1052389004, -1103483252, 1044014016, -1185623812, -1416839988, -1235231517, 1044000619, -1103483252, 1065353216, -1416839988, 1044000396, -1103483252, -1103483252, 1044065910, -1166022026, -1416839988, -1166610023, 1044063613, -1103483252, 1044085169, -1163554101, -1103483252, -1163615573, 1044084689, -1415753340, -1103483252, -1103483252, 1044000396, -1530674563, -1416839988, -1599121223, 1044000396, -1103483252, -1416839988, 1044000396, 0, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, 1065353216, -1416839988, 1044000396, -1103483252, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1758358451, -1416839988, -1103483252, -1847937581, 1044000396, -1263617743, 1044045727, -1171194459, -1103483252, -1103483252, -1416827918, -1171917758, 1044042880, -1416839988, 0, -1103483252, 1044000396, -1103483252, -1103483252, -1223220815, 924262833, -1103483252, -1764187712, 383295936, -1103483252, 1060777612, -1103483252, 1044138121, -1157202065, -1275395113, -1157045371, 1044140578, -1103483252, -1103483252, 1044000396, -2147479330, -1416839988, -2147483639, 1044000396, -1103483252, 1044068269, -1165717599, -1103483250, -1166038780, 1044065845, -1416838664, -1103483252, 1044004307, -1200325959, -1103483252, -1196709240, 1044005889, -1416839988, -1103483252, 1065353216, -1103483252, 1044000396, 0, 1052389037, -1103483252, -1103483252, 1065353216, -1103483252, 1044089117, -1163048779, -1103483252, -1416839988, -1163406415, 1044086323, -1416839988, 0, -1103483252, 1044000396, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, 0, -1416839988, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1065913784, 0, 1082231448, -1103483252, -1103483252, -1103483252, 0, -1223714092, 923769556, 0, -1103483252, 1057727209, -1103481510, 936997367, -1103483252, -1416735470, 1057727209, -1103481033, 940227016, 1065353216, 1082612749, -1103483252, -1416839988, -1103483252, -1416839988, -1416839988, -1065913784, 1065353216, -1103483252, -1103483252, 935703727, -1211779921, 0, 0, 1052389004, -1285321189, 1044035509, -1173805546, -1103483252, -1416839988, -1175250717, 1044031512, -1103483252, -1103483252, 1044014162, -1185474393, -1416839988, -1234870612, 1044000625, -1103483252, -1416839988, 1044000396, -1620082383, -1103483252, -1416839988, -1548531079, 1044000396, -1103483252, -1103483252, 1044039954, -1172666825, -1290019753, -1171708464, 1044043700, -1103483252, -1103483252, 1044000916, -1224601241, -1290021340, -1188992776, 1044010728, -1103483252, 1065353216, -1103483252, 1044000396, -1979545559, -1416839988, -1910762307, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1893079555, -1416839988, -1103483252, -1948581380, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 956354024, -1191129624, 236687925, -1910795723, 0, 0, 1065353216, -1416839988, 1044000396, -2008075180, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044031507, -1175253255, -1103483252, -1281025927, -1103483252, -1173810508, 1044035491, -1416839988, -2079680499, -1103483252, 1044000396, 912941841, -1234541807, -2147480921, 2727, -1103483252, -1103483252, -1103483252, -1222130260, 1057727376, -1103483252, -1103483252, -1208514517, 938969131, -1200800910, 946682738, -2008110660, 139372988, 1052389004, -1103483252, 973139123, -1174344525, -1188573690, 958909958, -1103483252, -1103483252, -1103483252, -1103483252, 1063828015, -1103483252, -1103483252, -1872438913, 275044735, 942857114, -1204626534, -1103483252, 940199323, -1207284325, -1899128880, 248354768, 1057727209, -1103483252, -1103483252, -1103483252, -1222130260, 1057727376, 968049308, -1179434340, -1235016322, 912467326, -1235011771, 912471877, 901256170, -1246227478, 1065353216, -1329848228, 817635420, -1103483252, -1188459947, 959023701, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, 907786183, -1239697465, -1232529692, 914953956, -1533990156, 613493492, 0, 0, 598921912, -1548561736, 946678329, -1200805319, 1052389004, -1103483252, 722938885, -1103483252, 808594238, 953680002, -1187980266, -1416839988, -1103490083, -1178624661, -1208904677, 938577872, -1103483252, -1416839988, -1103483896, -1222228421, 888837432, -1252742962, -1103483046, 911086376, 1070694194, -1416839988, -1103483252, -1416839988, -1218920922, 928204891, -1103485466, -1207247679, -1236698303, 910552324, -1103483252, -1416839988, -1416839988, -1416839988, 909677432, -1237468096, 1065353216, -1103483257, -1281712406, -1103483196, 895633847, -1103483196, 895638408, -1103485206, -1208549607, -1416839988, -1103483252, 831098405, 1075267027, -1103480595, 942018058, -1416839988, -1103481560, 936610497, -1103483252, -1416840188, -1416839988, -1416839988, -1103483252, -1416839988, -1103480566, 942138204, -1416839988, -1416839988, -1103484783, -1212176933, -1103484819, -1211884107, -1103483252, -1416839988, -1416839988, -1416839988, 1065353216, 1044000396, -1505008528, -1103483252, -1449237878, 1044000396, -1103483252, -1416839988, 1044044504, -1171501986, -1103483252, -1190771965, 1044008988, -1103483252, -1416839988, 1044094251, -1103483252, -1162391682, 1065353216, -1103483252, 1044000396, -1416839988, 1044000396, -1103483252, -1103483252, 1052389004, -1103483252, -1416839988, -1103483252, 1044000396, -1658426283, -1416839988, -1601137134, 1044000396, -1103483252, -1103486213, 1052395563, -1103483252, -1416839988, -1416839988, -1416839988, 1065353216, -1183106969, -1161334626, -1186138307, 1044115627, -1103483252, 1044000396, -1869818724, -1103483252, -1938774895, 1044000396, -1416839988, -1103483252, 1044001338, -1217690168, -1103483252, -1177285626, 1046329203, -1123255420, -1103483252, 1065353216, -1103483252, 1044066430, -1165952755, -1230400188, -1165643848, 1044069182, -1103483252, 950374310, -1103483252, -1197109338, -1869849526, 277634122, -1103483252, -1103483252, 1057727209, -1103483252, -1416839988, -1103486784, -1123241295, 1058302710, -1103484984, -1207866532, 1065353216, -1103483252, -1103483252, 925528851, -1221954797, 1052389004, 0, 0, 430071701, -1717411947, -1211914261, 935569387, -1222755507, 924728141, -1221940380, 925543268, 0, 0, -1103483252, -1103483252, 1052389004, 1065353216, -1103483252, 1044044739, -1171441822, -1413083928, -1171438822, 1044044751, -1103483252, 1065353216, -1103483252, 1044000396, -1399077823, -1416839988, -1449636145, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -2011630501, -1103483252, -1103483252, -1954883283, 1044000396, -1416839988, -1103483252, 1044056864, -1168337910, -1416839987, -1166755200, 1044063046, -1381374197, -1103483252, 1044000396, -1475934026, -1103483252, -1527376108, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044044637, -1171467962, -1103483252, -1416839988, -1174179651, 1044034044, -1103483252, -1416839988, 1044000396, -1309734341, -1087044365, -1253301646, 1063489699, -1103483252, 1044025699, -1178227036, -1103483252, -1178584893, 1044025000, -1416827342, -1103483252, 1065353216, -1103483252, 1044031431, -1175292153, -1111792847, -1171144808, 1049381106, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1318703601, -1243703727, -1103483252, -1260780988, 1044000534, -1087044365, -1103483252, 1063489686, -1335209259, -1416839988, -1406398372, 1044000396, -1103483252, -1103483252, -1193230454, 954253194, -1103483252, 884344627, -1263139021, 1052389004, 947097936, -1200385712, -1103483252, -1103483252, -1337823413, 809660235, 1052389004, -1103483252, 1044000598, -1236668172, -1343313275, -1174539407, 1044032901, -1103483252, -1103483252, 1044043887, -1171659958, -1416839988, -1173729636, 1044035802, -1103483252, 1044000396, -1331547014, -1103483252, -1389651105, 1044000396, -1416839988, -1103483252, 1044023690, -1179255563, -1103483252, -1187556888, 1044012128, -1416839988, -1103483252, -1103483252, -1103483252, -1336339461, 811144187, -1191436182, 956047466, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044035183, -1173888111, -1416839988, -1103483252, -1181643405, 1044019026, -1339581008, -1103483252, 1044040142, -1172618566, -1416839988, -1182504055, 1044017345, -1103483252, 1044124061, -1158575979, -1103483252, -1158077924, 1044128056, -1244696309, -1103483252, 1044000396, 0, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1065353216, -1103483252, 1044044739, -1171441764, -1413096080, -1171438888, 1044044750, -1103483252, 1065353216, -1103483252, 1044000396, -1399193761, -1416839988, -1449752765, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, 1044030130, -1175958323, -1103483252, -1103483252, -1178872183, 1044024439, -1416839988, -1103483252, 1044000396, -1788921392, -1416839988, -1836752579, 1044000396, -1416839988, -1103483252, 1044052944, -1169341275, -1103483252, -1169337086, 1044052961, -1412343840, -1103483252, 1044000396, 0, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044000396, -1377724170, -1103483252, -1330269802, -1323264689, 1044000396, -1103483252, -1331164654, 1044001153, -1220713598, -1416839988, -1308397914, 1044000396, -1103483252, 1044000396, -1735007974, -1103483252, -1803843168, 1044000396, -1103483252, -1416839988, 1044043258, -1171821079, -1103483252, -1171478372, 1044127134, -1163840293, -1103483252, 1052389004, -1103483252, -1103483252, 1044035506, -1173805537, -1103483252, -1103483252, -1172418321, 1044040957, -1258074545, -1103483252, 1082231448, -1343626057, -1065913784, -1405248629, 1044000396, -1416839988, -1103483252, -1103483252, 819640886, -1327842762, -1103483252, 944636270, -1202847378, 1052389004, -1789194554, 358289094, -1103483252, -1103483252, -1346199762, 801283886, 1052389004, -1103483252, 1044116251, -1159575683, -1416839988, -1159639054, 1044115756, -1103483252, 1065353216, -1103483252, 1044000396, -1416839988, 1044000396, -1103483252, 1044011274, -1188431724, -1103483252, -1251518410, 1044000453, -1416839988, -1103483252, 1044000396, -1419525545, -1103483252, -1355357914, 1046827227, -1121154753, -1103483252, -1103483252, -1103483252, -1192783567, 954700081, 789967737, -1357515911, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1618417733, -1299982791, -1103483252, -1559098535, 1044000397, -1300001763, -1103483252, 1044065076, -1166235768, -1416839420, -1166817377, 1044062803, -1103483252, 1044000396, -1314164084, -1103483252, -1361030794, 1044000396, -1416839988, -1103483252, 1044049173, -1170306794, -1103483252, -1168645904, 1046493731, -1122709796, -1103483252, 1065353216, -1103483252, 1044044740, -1171441637, -1413123425, -1171438951, 1044044750, -1103483252, 1044000396, -1399074943, -1103483252, -1449633330, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1519342706, -1103483252, -1103483252, -1458823953, 1044003349, -1204250783, -1103483252, 1044006494, -1195470196, -1416837168, -1180013119, 1044022216, -1281144467, -1103483252, 1044000396, -1885787215, -1103483252, -1822109256, 1044000396, -1416839988, -1103483252, 1044000396, -1534952842, -1103483252, -1476659307, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044000396, -1524965332, -1103483252, -1416839988, -1465184683, 1044000396, -1103483252, -1416837169, 1044000397, -1293292252, -1281149682, -1237892928, 1044000584, -1103483252, 1044026094, -1178024978, -1103483252, -1182649007, 1044017062, -1416839988, -1103483252, 1065353216, -1103483252, 1044024025, -1179084159, -1416839988, -1193142117, 1044007631, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044006074, -1196329725, -1305863818, -1103483252, -1174489373, 1044033000, -1305860139, -1103483252, 1044034737, -1174002393, -1416839988, -1207865672, 1044002467, -1103483252, -1103483252, 682219669, -1465263979, -1103483252, 967150691, -1180332957, 1052389004, 960026376, -1187457272, -1103483252, -1103483252, -1177595501, 969888147, 1052389004, 1052389004, -1103483252, -1103483252, 1044000660, -1232848945, -1103483252, -1103483252, -1177771946, 1044457802, -1143829044, -1103483252, 1044447672, -1176868830, -1144209646, -1205169871, 1044003125, -1416839988, -1103483252, 1044000396, -2147481964, -1103483252, -2147349295, 1044000396, -1416839988, -1103483252, 1044000396, -2133143397, -1103483252, -2147364594, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044001180, -1220277198, -1103483252, -1416839988, -1174551444, 1044032878, -1103483252, -1416839988, 1044000396, -1440019986, -1416839988, -1499229208, 1044000396, -1103483252, 1044020214, -1181035359, -1103483252, -1181309514, 1044019678, -1416674867, -1103483252, 1065353216, -1103483252, 1044021283, -1180488254, -1416839988, -1189803874, 1044009934, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044026505, -1177814551, -1416839988, -1103483252, -1215399284, 1044001535, -1416611355, -1103483252, 1044000397, -1297183301, -1416839988, -1363659491, 1044000396, -1103483252, -1103483252, 968438759, -1179044889, -1103483252, -1181096170, 966387478, 1052389004, -1179132043, 968351605, -1103483252, -1103483252, -1299536934, 847946714, 1052389004, -1103483252, 1044000396, -1305621741, -1416839988, -1364089261, 1044000396, -1103483252, -1103483252, 1044019792, -1181251468, -1416839988, -1231009675, 1044000716, -1103483252, 1044000396, -1318187687, -1103483252, -1376311667, 1044000396, -1103483252, -1416839988, 1044024958, -1178606302, -1103483252, -1177244167, 1044027619, -1342141306, -1103483252, -1103483252, -1103483252, -1323598571, 823885077, 935731696, -1211751952, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044028566, -1176758972, -1416839988, -1103483252, -1208218453, 1044002412, -1416839988, -1103483252, 1044000397, -1297778384, -1416839988, -1103483252, -1357475407, 1044000396, 1044081385, -1164038521, -1103483252, -1165939480, 1044066533, -1416839988, -1103483252, -1103483252, 1044000396, -1399947416, -1416839988, -1466678265, 1044000396, -1103483252, 1065353216, -1103483252, 1044044739, -1171441805, -1413091160, -1171438847, 1044044751, -1103483252, 1065353216, -1103483252, 1044000396, -1399077958, -1416839988, -1449636285, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1580071027, -1103483252, -1103483252, -1522700918, 1044000396, -1416839988, -1103483252, -1416839988, -1608189046, 1044000396, -1416839988, 1044000396, -1666500636, -1103483252, -1103483252, 1044200690, -1153197699, -1123496756, -1137417907, 1046980563, -1103483252, -1103483252, 1044000541, -1240369252, -1416839988, -1180795190, 1044020683, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044000410, -1268838574, -1075864298, -1103483252, -1197964685, 1073145162, -1167829570, -1103483252, 1044114723, -1168490003, -1416839988, -1169117039, 1044053820, -1103483252, 1044038863, -1172945980, -1103483252, -1174922971, 1044032152, -1416839988, -1103483252, 1065353216, -1103483252, 1044020448, -1180915307, -1416839988, -1213214924, 1044001802, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044062353, -1166932524, -1334681888, -1103483252, -1166349761, 1044064630, -1334659967, -1103483252, 1044030853, -1175587965, -1416839988, -1215510167, 1044001522, -1103483252, -1103483252, 946124934, -1201358714, -1103483252, 924383397, -1223100251, 1052389004, 539206937, -1103483252, -1608276711, -1103483252, -1178910266, 968573382, 1052389004, -1103483252, 1044000396, -1859696838, -1416839988, -1934099873, 1044000396, -1103483252, -1103483252, 1044071344, -1165323670, -1326917061, -1164850508, 1044075041, -1103483252, 1044024343, -1178921355, -1103483252, -1204505305, 1044003287, -1416839988, -1103483252, 1044000396, -1336805872, -1103483252, -1402739100, 1044000396, -1416839988, -1103483252, -1103483252, -1103483252, -1181977385, 965506263, -1339579668, 807903980, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044057266, -1168234794, -1416839988, -1103483252, -1170469623, 1044048537, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 1045065843, -1132327109, -1103483252, -1124827560, 1046116820, -1159872891, -1103483252, 1044024794, -1178690546, -1103483252, -1186658993, 1044013005, -1416839988, -1103483252, 1065353216, -1103483252, 1044044739, -1171441701, -1413103363, -1171438936, 1044044750, -1103483252, 1065353216, -1103483252, 1044000396, -1399048728, -1416839988, -1449607249, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, 0, -1103483252, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000396, -1445829240, -1416839988, -1507868121, 1044000396, -1416839988, -1103483252, 1044000396, -1412602812, -1103483252, -1463117235, 1044000396, -1416839988, -1103483252, 1044025127, -1178519862, -1103483252, -1178518367, 1044025130, -1103483252, -1413197351, 1052389004, -1103483252, -1103483252, 1044000396, -1436007945, -1103483252, -1103483252, -1376915681, 1044000396, -1327788927, -1103483252, 1044062471, -1166902424, -1416839936, -1166319917, 1044064747, -1329426831, -1103483252, 1065353216, -1103483252, 1044000396, -1394014163, -1416839988, -1444527376, 1044000396, -1103483252, 1044024858, -1178657793, -1103483252, -1178657810, 1044024858, -1103483252, -1413274769, 1052389004, -1103483252, -1103483252, -1103483252, 1044069819, -1165518989, -1413583859, -1103483252, -1165522710, 1044069789, -1413584779, -1103483252, 1044000396, -1303516814, -1416839988, -1376742089, 1044000396, -1103483252, -1103483252, -1103483252, 767297143, -1380186505, -1266029358, 881454290, 1052389004, -1447450089, 700033559, 924363097, -1223120551, -1103483252, -1103483252, 1052389004, -1103483252, 1044119745, -1159128457, -1416839988, -1159201866, 1044119171, -1103483252, 1065353216, -1103483252, 1044000396, -1416839988, 1044000396, -1103483252, 1044000397, -1297215079, -1103483252, -1240543364, 1044000539, -1334321185, -1103483252, 1044025045, -1178561704, -1103483252, -1213527492, 1044001764, -1416839988, -1103483252, -1103483252, -1103483252, 902249046, -1245234602, -1181915803, 965567845, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044035386, -1173836201, -1146307774, -1103483252, -1162343094, 1044448384, -1335185644, -1103483252, 1044081611, -1164009507, -1416839956, -1164340963, 1044079022, -1103483252, 1044000396, -1383969952, -1103483252, -1326089396, 1044000396, -1383522666, -1103483252, 1044044303, -1171553508, -1103483252, -1199562335, 1044004496, -1416839988, -1103483252, 1065353216, -1103483252, 1044044739, -1171441803, -1413091293, -1171438847, 1044044751, -1103483252, 1065353216, 1065353216, -1103483252, 1044000396, -1399077947, -1416839988, -1449636276, 1044000396, -1103483252, -1103483252, 1044032604, -1174691442, -1416839988, -1237687230, 1044000582, -1103483252, -1103483252, 1044001593, -1214924277, -1324887415, -1173525602, 1044036599, -1103483252, 1044000396, -1533891030, -1103483252, -1602052645, 1044000396, -1416839988, -1103483252, 1044000396, -2147483647, -1103483252, -2147483646, 1044000396, -1408382282, -1103483252, 1065353216, 1065353216, -1103483252, 1044043842, -1171671546, -1408395442, -1171616121, 1044044058, -1103483252, 1044108482, -1160570047, -1103483252, -1160417007, 1044109678, -1397439203, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044125746, -1158360237, -1103483252, -1416835960, -1158626214, 1044123668, -1103483252, -1416835957, 1044000396, -1455378359, -1416839988, -1506552583, 1044000396, -1103483252, -1103483778, -1224515757, 1052389004, -1103482070, 932436892, -1416711039, -1416964906, 1065353216, -1537636249, 609847399, -1103483252, -1103483252, 925337888, -1222145760, -1103483252, 1057727209, -1103483252, -1416840138, -1103483252, -1408382282, 1057727209, -1103483347, -1245904774, 1065353216, -1103483252, -1103483252, 1, -2147483647, -1218460332, 929023316, 1052389004, -1416839955, 1044047603, -1170708557, -1103483252, -1334319761, -1170766974, 1044047375, -1103483252, -1416839988, 1044000396, 0, -1103483252, -1416839988, 0, 1044000396, -1103483252, -1416499543, 1044017500, -1182424895, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044000542, -1240335397, -1103483252, -1217881146, -1103483252, -1185736418, 1044014836, -1416839988, -1214695089, -1103483252, 1044001621, -1103483252, 1044039655, -1172743351, -1338534002, -1171770370, 1044043456, -1103483252, -1103483252, 1044039508, -1172780869, -1361165081, -1171799828, 1044043341, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1478544141, -1416839988, -1103483252, -1537301144, 1044000396, -1416839988, -1103483252, 1044000396, -1809475920, -1416839988, -1761627464, 1044000396, -1103483252, -1103483252, 1044000481, -1247065331, -1416839988, -1308560344, 1044000396, -1103483252, 1065353216, -1103483252, 1044003367, -1204176166, -1224217022, -1175138589, 1044032275, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1354278610, -1416839988, -1103483252, -1406440300, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 385516965, -1761966683, -1249345361, 898138287, 968378564, -1179105084, 0, 0, 1065353216, -1416839988, 1044000396, 0, -1103483252, -1416839988, 0, 1044000396, -1103483252, -1416839988, 1044001723, -1213861017, -1103483252, -1096276143, -1183166998, 1057140464, -1103483252, -1103483252, 1044085171, -1163553878, -1415751633, -1163615269, 1044084691, -1103483252, -1103483252, 1044000396, -1530694092, -1416839988, -1599138824, 1044000396, -1103483252, -1416839988, 1044000396, 0, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1335750754, 1044047374, -1170767171, -1103483252, -1416839958, -1103483252, -1170708728, 1044047603, -1416839988, 0, -1103483252, 1044000396, -1103483252, 1044000396, -1513371864, -1416839988, -1582200174, 1044000396, -1103483252, -1103483252, 1044000396, 0, -1134796792, 0, 1044903052, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044109901, -1160388474, -1400701303, -1103483252, -1160257634, 1044110923, -1400451458, -1103483252, 1044089266, -1163029682, -1256754235, -1162128861, 1044096342, -1103483252, -1103483252, 1044000528, -1241245593, -1416839988, -1308028310, 1044000396, -1103483252, 1065353216, -1103483252, 1044002888, -1206141109, -1132191752, -1178501324, 1045107530, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044132735, -1157546774, -1342176652, -1103483252, -1157471840, 1044133906, -1343487166, -1103483252, 1044059415, -1167684850, -1416839988, -1184483858, 1044015129, -1103483252, 949008697, -1198474951, -1244477805, 903005843, 966079731, -1181403917, -1174009266, 973474382, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, 0, 0, 914418904, -1233064744, 1063828015, -1103483252, -1103483252, -1103483252, -1103483252, -1516784429, 630699219, 923756123, -1223727525, 1060777612, -1103483252, -1103483252, 940205808, -1207277840, -1357375966, 790107682, -1103483252, -1103483252, 1060777612, 0, 0, -1187093704, 960389944, 0, 0, -1103483252, -1103483252, 908503184, -1238980464, 1052389004, -1180168428, 967315220, 971093984, -1176389664, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1238980445, 908503203, 958888076, -1188595572, 960671629, -1186812019, -1232541703, 914941945, -1534004681, 613478967, 0, 0, 1052389004, 815960446, -1331523202, -1175399875, 972083773, 940202559, -1207281089, -1483869116, 663614532, -1103483252, -1103483252, -1103483252, 1057727209, -1103483294, -1255696722, -1103483252, -1339684299, 1070691542, -1103483252, 722945309, -1103472742, 958675812, -1250549100, 896918665, 941974154, -1201698436, -1103483252, -1416860343, -1416839988, -1416839988, -1103483252, 774762369, -1416839988, -1416839988, -1416839988, -1416839988, -1103483047, 911068699, 896946106, -1250523056, -1103483701, -1226814586, 940992572, -1206335988, -1103484165, -1218166497, -1189360338, 958123281, 1065353216, -1103478070, 950138176, -1103474271, 957110053, 1076768638, -1103483257, -1281196288, -1103489366, -1195438084, -1416839988, -1416839988, -1201218434, 946265214, -1103484839, -1211735131, -1103484870, -1211484053, -1103483235, 881271221, -1103488028, -1197066027, 940277697, -1096275027, -1103483252, -1416840187, -1416839988, -1416839988, -1103483252, -1416840810, -1103483252, -1134796792, -1103483226, 886136883, -1103486430, -1132166335, 1065353216, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, 0, 0, -1417430499, 730053149, 852719013, -1294764635, 966801954, -1180681694, -1103483252, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 918634338, -1228849310, -1103483252, 1060777612, -1103483254, -1297995436, -1103483252, -1327739679, 936384698, -1211098171, -1103483252, 795517729, 1063916453, -1103483252, -1416839988, -1103521988, -1145068248, -1207789343, 939694070, 1065353216, -1399472928, 748010720, -1348682702, 798800946, -1308270470, 839213178, -1225129740, 922353908, 905183381, -1242300267, -1459559875, 687923773, 1065353216, -1103483252, -1416839988, -1416743797, -1416936179, -1103483252, -1425245668, 1063828015, -1103483252, 733088822, -1103483241, 876435151, -1315951295, 831527054, -1103482292, 930087027, 1065353216, -1103483252, 1044032607, -1174690224, -1416839988, -1237685227, 1044000582, -1103483252, -1103483252, 1044001598, -1214890102, -1273477626, -1173644597, 1044036144, -1103483252, 1044000396, -1526094604, -1103483252, -1594406673, 1044000396, -1416839988, -1103483252, 1044044262, -1171563884, -1103483252, -1171566978, 1044044250, -1413460803, -1103483252, 1065353216, -1103483252, 1044000396, 0, -1413461410, 0, 1044000396, -1103483252, 1044109495, -1160440370, -1103483252, -1160498313, 1044109043, -1415341660, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044129817, -1157839192, -1103483252, -1336753704, -1157797271, 1044130145, -1103483252, -1334842744, 1044000396, -1349338782, -1416839988, -1398258369, 1044000396, -1103483252, -1103483049, 910890331, 1052389004, -1103483747, -1225303145, -1333555800, 783766355, 1065353216, -1530100389, 617383259, -1103483252, -1103483252, -1233544890, 913938758, -1103483252, 1057727209, -1103483252, -1416840267, -1103483247, 866874734, 1057727209, -1103483252, -1413461410, 1065353216, -1103483252, -1103483252, 0, 0, -1238947532, 908536116, 1052389004, -1416839988, 1044031515, -1175249377, -1103483252, -1287595214, -1173803261, 1044035518, -1103483252, -1416839988, 1044000396, -1621802754, -1103483252, -1416839988, -1549818927, 1044000396, -1103483252, -1344562578, 1044019832, -1181230724, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839666, 1044000399, -1284466017, -1103483252, -1307228890, -1103483252, -1227521050, 1044000823, -1416839988, -1214994299, -1103483252, 1044001585, -1103483252, 1044033177, -1174401768, -1416839988, -1183393057, 1044016194, -1103483252, -1103483252, 1044013999, -1185641393, -1416839988, -1235273526, 1044000619, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1825288961, -1416839988, -1103483252, -1777650389, 1044000396, -1416839988, -1103483252, 1044000396, -1638015592, -1416839988, -1590997861, 1044000396, -1103483252, -1103483252, 1044000482, -1247004333, -1416839988, -1308512659, 1044000396, -1103483252, 1065353216, -1103483252, 1044000602, -1236362171, -1416839988, -1305867893, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044001091, -1221733259, -1204775779, -1103483252, -1172292692, 1044044241, -1333029734, -1103483252, 1044122494, -1158776511, -1416839950, -1159325669, 1044118204, -1103483252, 556258596, -1591225052, -1249296269, 898187379, -1239095077, 908388571, -1211017491, 936466157, 1065353216, -1416839985, 1044000397, -1293260556, -1103483252, -1364807198, -1236759374, 1044000596, -1103483252, -1344562578, 1044020364, -1180958422, -1103483252, -1416839988, -1214260312, 1044001675, -1103483252, -1103483252, 1044085165, -1163554628, -1415762634, -1163616542, 1044084681, -1103483252, -1103483252, 1044000396, -1530668215, -1416839988, -1599115478, 1044000396, -1103483252, -1416839988, 1044000396, -1550819426, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1286949161, 1044035515, -1173803945, -1103483252, -1416839988, -1103483252, -1175249762, 1044031514, -1416839988, -1623139265, -1103483252, 1044000396, -1103483252, 1044000638, -1234001785, -1416839988, -1192212574, 1044008085, -1103483252, -1103483252, 1044043038, -1171877217, -1264447068, -1167216849, 1044061263, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044009067, -1190691062, -1223307619, -1103483252, -1169907101, 1044051333, -1416839522, -1103483252, 1044139267, -1157128761, -1302878826, -1156999253, 1044141291, -1103483252, -1103483252, 1044000508, -1243503567, -1416839988, -1308389767, 1044000396, -1103483252, 1065353216, -1103483252, 1044003394, -1204066654, -1264417341, -1174986743, 1044032048, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -2147483647, -1416839988, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, -1256377455, 891106193, -1246496868, 900986780, 968358337, -1179125311, 0, 0, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, 954860146, -1192623502, 0, 0, 1063828015, -1103483252, -1103483252, -1103483252, -1103483252, 954774173, -1192709475, 973896685, -1173586963, 1060777612, -1103483252, -1103483252, -1188587079, 958896569, 973163056, -1174320592, -1103483252, -1103483252, 1060777612, 597637424, -1549846224, -1184583275, 962900373, 906606013, -1240877635, -1103483252, -1103483252, -1200800009, 946683639, 1052389004, -1180167586, 967316062, 971125484, -1176358164, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, 946684104, -1200799544, 915907630, -1231576018, -1184228446, 963255202, -1232464963, 915018685, -1533985434, 613498214, -1550844112, 596639536, 1052389004, 1010133878, -1137349770, -1189988948, 957494700, -1187036281, 960447367, 369648631, -1777835017, -1103483252, -1103483252, -1103483252, 1057727209, -1103480175, 943740876, -1103677601, -1147775702, 1070706042, -1103483252, 723026275, -1103472741, 958676531, 910943916, -1236342243, 904919552, -1242487661, -1103483252, -1416839988, -1416839988, -1416839988, -1103490479, -1189278257, -1205634469, 941848900, 896796796, -1250685500, -1103483045, 911183093, -1236450409, 910825655, -1103488955, -1195053196, 939584946, -1207895252, -1103483252, -1416839988, -1416839988, -1416839988, 1065353216, -1103483252, 790930299, -1103480821, 941094016, 1075267029, -1103483257, -1281880847, -1103488836, -1196505366, -1416839988, -1416839988, -1201557066, 945926472, -1103478511, 949234674, -1103480599, 942003919, -1103483235, 881317356, -1103483211, 891561328, -1201164962, 946318576, -1103483252, -1416840188, -1416839988, -1416839988, -1103483252, -1411093240, -1103493969, -1188576751, -1103483230, 884118973, -1103488337, -1197504425, 1065353216, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, -1865689201, 281794447, 935509996, -1211973652, -1103483252, 1060777612, 624675194, -1522808454, 1004882815, -1142600833, -1205758816, 941724832, -1203914675, 943568973, -1103483252, -1103483252, 1052389004, 963335048, -1184148600, -1200896286, 946587362, -1184871575, 962612073, 0, 0, -1103483252, -1103483252, -1277728882, 869754766, -1354535560, 792948088, 1052389004, -1103479126, 947973947, 1063828015, -1103478961, 948313011, -1103484917, -1211100456, -1196976876, 950506650, -1103485391, -1207588058, -1103477558, 951185985, -1416839988, -1416839988, 1065353216, -1103483252, -1416839988, 1076637327, -1416839988, -1103552199, -1123220969, -1103488333, -1197553571, -1416839988, -1103484459, -1075864147, -1168168277, -1213898166, -1103483252, -1416839988, 1065353216, -1103483252, 1044099635, -1161702441, -1400541392, -1161537725, 1044100922, -1103483252, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 1044000396, -1340403636, -1103483252, -1409306842, 1044000396, -1416839988, -1103483252, 1044042313, -1172062968, -1103483252, -1172782388, 1044039502, -1416839969, -1103483252, 1065353216, -1103483252, 1044042680, -1171968838, -1416839970, -1172680161, 1044039902, -1103483252, 1044098169, -1161890142, -1103483252, -1161273748, 1044102985, -1345510973, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044000712, -1231142419, -1103483252, -1132361633, -1174211123, 1045095053, -1103483252, -1132405980, 1045125732, -1165477397, -1416839988, -1182424413, 1044017501, -1103483252, -1103485174, -1208996841, 1053447364, -1103489852, -1132308836, -1132319124, 959030335, 1065353216, -1343128302, 804355346, -1103483252, -1103483252, 942990219, -1204493429, -1103483252, 1057727209, -1103483252, 788934196, -1103482086, 932300074, 1057727209, -1103482088, 932288157, 1065353216, -1103483252, -1103483252, -1211515692, 935967956, 969925420, -1177558228, 1052389004, -1416839988, 1044000396, -1655457270, -1103483252, -1103483252, -1416839988, -1606375207, 1044000396, -1310230695, 1044013204, -1186455782, -1103483252, -1416839738, -1103483252, -1190040626, 1044009703, -1416839988, 1044000396, 0, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416838979, 1044047480, -1170740004, -1103483252, -1293299610, -1103483252, -1170797497, 1044047258, -1416839988, 0, -1103483252, 1044000396, -1103483252, 1044000396, -1480479005, -1416839988, -1423346662, 1044000396, -1103483252, -1103483252, 1044000396, -1400168682, -1070263986, -1335808143, 1077982263, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044088014, -1163190030, -1381712712, -1103483252, -1161868771, 1044098336, -1381714190, -1103483252, 1044047705, -1170682417, -1416839988, -1228876495, 1044000781, -1103483252, -1103483252, 1044000459, -1250097240, -1416839987, -1308025676, 1044000396, -1103483252, 1065353216, -1103483252, 1044002048, -1211197394, -1077172226, -1182155938, 1071838827, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1490585904, -1416839988, -1103483252, -1433161776, 1044000396, -1416839988, -1103483252, 1044000396, -1576116398, -1416839988, -1608281680, 1044000396, -1103483252, -1174000024, 973483624, -1253490294, 893993354, 962159606, -1185324042, -1576786393, 570697255, 1065353216, -1201152249, 1044400933, -1144929415, -1103483252, -1416839988, -1150257720, 1044246627, -1103483252, -1416839988, 1044000405, -1273206715, -1103483252, -1077047050, -1202136293, 1071962233, -1103483252, -1103483252, 1044085171, -1163553873, -1415751575, -1163615261, 1044084691, -1103483252, -1103483252, 1044000396, -1530694390, -1416839988, -1599139093, 1044000396, -1103483252, -1310230695, 1044008872, -1190891593, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044000396, 0, -1103483252, -1416839988, -1103483252, 0, 1044000396, -1416839738, -1200187490, -1103483252, 1044004341, -1103483252, 1044076368, -1164680712, -1416839988, -1164992852, 1044073929, -1103483252, -1103483252, 1044000396, -1792793717, -1312596763, -1732716428, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, 0, -1416839988, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000396, -1688744116, -1416839988, -1641293121, 1044000396, -1103483252, -1103483252, 1044000460, -1249879369, -1416839988, -1308001623, 1044000396, -1103483252, 1065353216, -1103483252, 1044000890, -1225317863, -1312596764, -1189086881, 1044010634, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044101800, -1161425298, -1328301733, -1103483252, -1160579158, 1044108411, -1328301756, -1103483252, 1044000396, 0, -1416839931, 0, 1044000396, -1103483252, 505081873, -1642401775, -1253297546, 894186102, 956195075, -1191288573, 0, 0, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, 411306825, -1736176823, 945843632, -1201640016, 1063828015, -1103483252, -1103483252, -1103483252, -1103483252, -1224970235, 922513413, 0, 0, 1060777612, -1103483252, -1103483252, 809224648, -1338259000, 714236108, -1433247540, -1103483252, -1103483252, 1060777612, -1205568233, 941915415, 0, 0, -1159888009, 987595639, -1103483252, -1103483252, 0, 0, 1052389004, 926891225, -1220592423, 0, 0, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, 540890489, -1606593159, -1238987933, 908495715, 943403754, -1204079894, -1232542103, 914941545, -1534004903, 613478745, -1201494616, 945989032, 1052389004, -1189962029, 957521619, -1403345323, 744138325, 722333725, -1425149923, 952320704, -1195162944, -1103483252, -1103483252, -1103483252, 1057727209, -1103483252, 815866047, -1103477785, 950721618, 1070691885, -1103483252, 722945280, -1103483774, -1224574600, -1416839988, -1416839988, -1251466335, 895538444, -1103487326, -1199661077, -1186695436, 960788210, -1103483252, -1416839983, -1416839988, -1416839988, -1172325457, 974208446, -1103483047, 911068105, -1416839988, -1416839988, -1103483252, -1416839988, -1416839988, -1416839988, -1103486272, -1203979376, -1328301756, -1416839931, 1065353216, -1103484328, -1215927166, 1090927846, -1103483252, -1448751549, -1103483257, -1281188504, -1103483252, -1416839988, -1218880177, 928596063, -1416839988, -1416839988, -1103483252, -1415987940, -1103483252, -1070263986, -1103483240, 877037158, -1103485316, -1077171968, 921198153, -1077046992, -1103483252, -1416840187, -1218305208, 929171032, -1103481319, 938587901, -1103483252, -1312596763, -1103483240, 877229044, -1103484856, -1211594084, 1065353216, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1310649287, 836834361, -1183868850, 963614798, -1103483252, 968728387, -1178755261, 144702, -2147338946, -1230240833, 917242815, -1180709208, 966774440, -1103483252, -1103483252, 1052389004, -2138861763, 8621885, -1442683113, 704800535, -1191734127, 955749521, -1299072710, 848410938, -1103483252, -1103483252, -1211268526, 936215122, -1172096651, 975386997, 1052389004, -1103483061, 910126617, 1063828015, -1103479826, 945169012, -1103477983, 950316204, -1316171854, 831307235, -1103479511, 946461013, -1103477553, 951195459, -1324046285, 823428356, 1065353216, -1103484908, -1143776048, -1144155526, 936601697, -1103483252, -1416839988, -1103483252, -1416839988, 1064040648, -1103491244, -1191591796, -1416517566, -1417162410, -1103483252, 829383951, 1065353216, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, -1103483252, 1044128413, -1158018944, -1416839988, -1158493140, 1044124708, -1103483252, 1044000396, -1675041789, -1103483252, -1625707721, 1044000396, -1416839988, -1103483252, 1044008760, -1191006263, -1103483252, -1241038980, 1044000531, -1416839988, -1103483252, -1103483252, -1103483252, 521602978, -1625880670, -1194527078, 952956570, 1052389004, 1052389004, -1103483252, -1103483252, -1103483252, 1044044003, -1171630354, -1412974101, -1103483252, -1171626076, 1044044019, -1413064258, -1103483252, 1044027098, -1177510852, -1416839988, -1103483252, -1223007579, 1044001013, 1044044739, -1171441801, -1103483252, -1171438842, 1044044751, -1413091084, -1103483252, 1065353216, -1103483252, 1044000396, -1399075617, -1416839988, -1449633898, 1044000396, -1103483252, -1103483252, 1044001112, -1221394479, -1313762305, -1170885030, 1044046914, -1103483252, 1044018809, -1181754454, -1103483252, -1231501602, 1044000701, -1416839988, -1103483252, -1103483252, 1044102253, -1161367415, -1416839982, -1162564812, 1044092898, -1103483252, 1044000396, -1320913300, -1103483252, -1392161099, 1044000396, -1103483252, -1416839988, 1044000396, 0, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044048006, -1170605515, -1103483252, -1169774322, 1044051253, -1343514181, -1103483252, 1065353216, -1103483252, 1044004482, -1199609405, -1085337029, -1172791191, 1065206790, -1103483252, 1044122108, -1158825998, -1103483252, -1158358494, 1065062460, -1085502932, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044098446, -1161854664, -1103483252, -1416839988, -1163125588, 1044088517, -1103483252, -1416839988, 1044000396, -1455442418, -1416839988, -1519370568, 1044000396, -1103483252, -1103488207, -1085501694, 1066717369, -1103479150, 947926340, -1416787685, -1416892291, 1065353216, 0, 0, -1103483252, -1103483252, -1214068695, 933414953, -1103483252, 1057727209, -1103483252, -1416839988, -1103484889, -1211325629, 1068325522, -1103488522, -1085335712, 1065353216, -1103483252, -1103483252, 971516062, -1175967586, -1196027021, 951456627, 1052389004, 1044000396, -1103483252, -1416839988, -1103483252, 1052389339, -1103483252, -1222130260, -1416839289, 1044038854, -1172948478, -1103483252, -1298019062, -1103483252, -1172990280, 1044038692, 1044001100, -1221584403, -1103483252, -1180942947, 1044020395, -1325260679, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1305253460, -1416839988, -1103483252, -1363709269, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 1044000875, -1225817869, -1103483252, -1189144346, 1044010578, -1325260679, -1103483252, 1065353216, -1416839988, 1044000396, -1103483252, -1416839988, 1044000396, -1103483252, -1103483252, 1044095312, -1162255770, -1416839988, -1162259126, 1044095286, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, 0, -1416839988, -1103483252, 0, 1044000396, -1416839984, -1103483252, 1044088733, -1163097979, -1358929213, -1161806966, 1044098819, -1103483252, -1103483252, 1044000444, -1254113569, -1416839987, -1311758632, 1044000396, -1103483252, 1065353216, -1103483252, 1044001084, -1221850805, -1416839988, -1182921337, 1044016655, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, 0, -1416839988, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000851, -1226577047, -1369222646, -1170707754, 1044047606, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044109568, -1160431095, -1085894597, -1103483252, -1160182255, 1064667233, -1416839608, -1103483252, 1044109795, -1160402049, -1305478203, -1160349241, 1044110208, -1103483252, -1416839988, 1044000396, -1103483252, 1065353216, -1103483252, 1044001821, -1213063576, -1416839988, -1291480514, 1044000398, -1103483252, -1416839605, 1044049855, -1170132251, -1103483252, -1305394293, -1170182583, 1044049659, -1103483252, -1416839988, 1044000396, -1675044641, -1103483252, -1416839988, -1625710316, 1044000396, -1103483252, -1103483252, 1044095235, -1162265632, -1416839988, -1162270007, 1044095201, -1103483252, -1085411535, 1062072116, -1272895283, -1416839988, -1351049374, 1044000396, -1103483252, -1416839925, 1044022169, -1180034586, -1103483252, -1326776628, -1178990858, 1044024207, -1103483252, -1103483252, 1044085171, -1163553837, -1415751351, -1163615214, 1044084692, -1103483252, -1103483252, 1044000396, -1530694521, -1416839988, -1599139231, 1044000396, -1103483252, -1416839988, 1044032675, -1174655501, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044000396, 0, -1103483252, -1416839988, -1103483252, 0, 1044000396, -1226994699, -1172661598, -1103483252, 1044040417, -1240432701, 907050947, 932197392, -1215286256, -1103483252, -1103483252, 0, 0, 1052389004, -1213687886, 933795762, -1103483252, -1274533271, 872950377, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, -1222130260, 1057727376, 0, 0, -1103483252, -1103483252, -1103483252, -1103483252, -1267676450, 879807198, -1103483252, 1063828015, 952167906, -1195315742, -1256681843, 890801805, 961718313, -1185765335, 974110052, -1173373596, 1065353216, 0, 0, 956064084, -1191419564, -1230035621, 917448027, -1215407213, 932076435, 1065353216, -1103483252, -1103483252, -1103483252, -1269984161, 877499487, 0, 0, -1103483252, 1060777612, -1196465742, 951017906, -1323491021, 823992627, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, 973771806, -1173711842, -1184671639, 962812009, 964246091, -1183237557, -1310167645, 837316003, -1103483252, -1103483252, -1103483252, 1057727209, -1103483252, -1103483252, -1242359684, 905123964, 521600428, -1625883220, -1232543718, 914939930, -1534005000, 613478648, 943382890, -1204100758, 1052389004, -1103483252, -1416839988, 1075469886, -1103483252, 722951764, -1103493579, -1188996524, -1103479510, 946464562, -1255736931, 891415331, -1103483252, 829881916, -1416839988, -1416839988, -1103483252, -1416839988, 947160274, -1200323341, -1103483252, -1416839988, 958109293, -1189374351, -1103486545, -1085893773, 926856905, -1220615479, -1253019482, 894282630, -1416839988, -1416839988, -1103483047, 911065741, -1416839988, -1416839988, 1065353216, -1103481582, 936426481, -1103483257, -1281184218, -1103479694, 945709773, -1103483252, 807074123, -1416839988, -1103486596, -1202651317, -1103484879, -1211406924, 1077878481, -1416839988, -1416839988, -1103483239, 878048866, -1103483243, 873873354, -1103485342, -1207790807, -1416839988, -1103482968, 915275820, -1103483233, 882444749, -1085411535, 851836843, 928856534, -1218625233, -1103483252, -1416840187, 948350094, -1198226098, 1065353216, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, 1060777612, 0, 0, -1225421429, 922062219, -1103483252, 683605572, -1463878076, 325295969, -1822187679, -1196555294, 950928354, 872965137, -1274518511, -1103483252, -1103483252, 1052389004, 667225496, -1480258152, 906151751, -1241331897, -1187844155, 959639493, -1103483252, -1103483252, -1180559906, 966923742, 935934149, -1211549499, -1457177609, 690306039, 1052389004, -1103479790, 945319197, 1063828015, -1103478310, 949645791, -1103488987, -1196213682, -1196216094, 951266192, -1103480039, 944298173, -1103483261, -1274873753, -1197028063, 950455585, 1065353216, -1103483252, -1204250783, 947055825, -1200406922, -1103483252, -1416839988, -1103483252, -1416826452, 1063828755, -1103483252, -1416839988, 894080620, -1252066017, -1103483252, -1416839988, 1065353216, 1044141764, -1156968950, -1103483252, -1156904744, 1044142767, -1103483252, -1350185179, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 1044000396, 0, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044043034, -1171878410, -1103483252, -1173923251, 1044035046, -1416839988, -1103483252, 1065353216, -1103483252, 1044039929, -1172673132, -1416839988, -1173894135, 1044035160, -1103483252, 1044076650, -1164644532, -1103483252, -1163019729, 1047054450, -1120601656, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044000397, -1302025625, -1103483252, -1097489210, -1247175775, 1056095287, -1103483252, -1097701716, 1055882738, -1342420073, -1416839988, -1392992980, 1044000396, -1103483252, -1103486922, -1120586976, 1065118875, -1103483272, -1097489200, -1097701716, 788877479, 1065353216, 0, 0, -1103483252, -1103483252, 957153061, -1190330587, -1103483252, 1057727209, -1103483252, -1416839988, -1103479983, 944524913, 1057727209, -1103481420, 937759948, 1065353216, -1103483252, -1103483252, -1204318649, 943164999, 897619480, -1249864168, 1052389004, 1044011756, -1187938610, -1301132719, -1103483252, -1225090242, 1044000897, -1416839988, -1103483252, -1416839988, 1044000667, -1232635921, -1103483252, -1416839988, -1188501743, 1044011205, -1103483252, -1416839510, 1044044300, -1171554253, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, 1044000396, 0, -1416839988, -1103483252, -1103483252, 0, 1044000396, -1416839988, -1302507573, -1171552161, -1103483252, 1044044309, -1103483252, 1044009008, -1190751422, -1105372577, -1172169994, 1051465091, -1103483252, -1103483252, 1044000420, -1262454933, -1416839988, -1204379719, 1044003318, -1103483252, 1052389004, -1103483252, -1103483252, 1044000396, -1458384245, -1103483252, -1103483252, -1398097422, 1044000396, -1416839988, -1103483252, 1045150033, -1131653592, -1416839988, -1144133196, 1044422105, -1416839988, -1103483252, -1103483252, 1044003093, -1205299331, -1105318762, -1173919881, 1051488580, -1103483252, 1065353216, -1103483252, 1044031639, -1175185762, -1416839988, -1218375300, 1044001296, -1103483252, 1052389004, -1103483252, -1103483252, 1044001089, -1221761015, -1103483252, -1103483252, -1172073682, 1044042380, -1243918225, -1103483252, 1044089555, -1162992757, -1416839895, -1161906525, 1044098041, -1322550583, -1103483252, -1141270143, 1006213505, 970141060, -1177342588, -1178856967, 968626681, 950082087, -1197401561, 1065353216, -1065913784, 1082232154, -1179613894, -1103483252, -1416839988, -1206476963, 1044002806, -1103483252, 1044085179, -1163552898, -1103483252, -1163613671, 1044084704, -1415738678, -1103483252, -1103483252, 1044000396, -1530670206, -1416839988, -1599117555, 1044000396, -1103483252, -1416839988, 1044000396, -1623187843, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, 1044031530, -1175241536, -1416839988, -1103483252, -1103483252, -1173788742, 1044035572, -1299807825, -1416839988, -1550855796, -1103483252, 1044000396, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, -1103483252, 1044034446, -1174076868, -1416839988, -1182650760, 1044017059, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1416839895, 1044000396, -1103483252, -1103483252, 1044116675, -1159521387, -1103483252, -1416839988, -1159580431, 1044116214, -1103483252, -1283475058, 1044078460, -1164413430, -1416839988, -1169356555, 1044052885, -1103483252, -1103483252, 1044000517, -1242379034, -1416839988, -1308239887, 1044000396, -1103483252, 1065353216, -1103483252, 1044000482, -1247027978, -1416839988, -1308531507, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1322545643, 1044000396, -1103483252, -1103483245, 1044002064, -1211126593, -1416839988, -1103483252, -1264331334, 1044000416, -1416839988, -1103483252, 1044000396, -1558024034, -1416839988, -1500549240, 1044000396, -1103483252, -1181838951, 965644697, -1245597870, 901885778, -1249315488, 898168160, 646851239, -1500632409, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1186974669, 960508979, -1103483252, -1215178185, 932305463, 1063828015, -1103483252, -1103483252, -1103483252, 0, 0, -1103483252, 918017964, -1229465684, 1060777612, -1103483252, -1103483252, 943005385, -1204478263, 973178972, -1174304676, -1103483252, -1103483252, 1060777612, 956833384, -1190650264, 865677978, -1281805670, -1103483252, -1103483252, 946694637, -1200789011, 1052389004, 908815348, -1238668300, 0, 0, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1182777534, 964706114, 0, 0, -1182225635, 965258013, -1232632409, 914851239, -1533986613, 613497035, 596603261, -1550880387, 1052389004, -1319448801, 828034847, 948128432, -1199355216, 969062309, -1178421339, 745746091, -1401737557, -1103483252, -1103483252, -1103483252, 1057727209, -1103479842, 945103501, -1103483252, 820642730, -1103483252, 722953557, -1103484084, -1219496795, 950903182, -1196578527, -1416839988, -1416839988, -1103483252, -1406773164, -1152144683, 995338965, -1103491274, -1191307566, 944778938, -1202704024, -1103483049, 910933664, 913488505, -1233926271, 1070691436, -1416839895, -1103482423, 927940051, -1192955249, 954520216, -1322545643, -1103482771, 921504961, -1416839988, -1416839988, 1065353216, -1103483252, -1121154753, -1103485539, -1122700650, 1087617780, -1103483257, -1282167970, -1103483252, -1416839988, 937715531, -1209768116, 861439889, -1282937265, -1103491215, -1105364615, -1103483252, -1392830379, -1103488188, -1105313827, -1103476982, 952365159, -1065913616, 942158217, -1103483252, -1416840188, -1416839988, -1416839988, -1103483252, -1416839988, -1103478166, 949940123, -1103483228, 885016427, -1103483235, 881300240, 1065353216, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, 918055721, -1229427927, -1103483252, 1060777612, -1199575218, 947908430, 875049774, -1272433874, -1739425427, 408058221, 584813021, -1562670627, -1103483252, -1103483252, 1052389004, 0, 0, -1224664130, 922819518, 930751726, -1216731922, -1223138502, 924345146, -1103483252, -1103483252, -1198295539, 949188109, -1347079150, 800404498, 1052389004, -1103483252, -1416839988, -1103483590, -1163797013, -1103485375, -1207519041, -1065913784, 781514326, 1083759230, -1103483252, -1416839988, -1103483252, -1299982791, -1211110300, 936364928, 1065353216, -1103481656, 935822756, -1416839988, -1416839988, -1103483258, -1279571016, -1103483252, -1416839988, 1063828015, -1103483252, -1324593714, -1234128730, 913349536, -1103482388, 928512816, 1065353216, -1103483252, 1044000399, -1287221531, -1416839988, -1344700738, 1044000396, -1103483252, -1103483252, 1044046837, -1170904852, -1416839988, -1178934533, 1044024317, -1103483252, 1044046394, -1171018209, -1103483252, -1178131587, 1044025885, -1416839988, -1103483252, 1044000396, -1524686808, -1103483252, -1454139438, 1044000396, -1416839988, -1103483252, 1065353216, -1103483251, 1044000397, -1327950639, -1416839988, -1393462652, 1044000396, -1103483252, 1044000400, -1283378349, -1103483252, -1341054134, 1044000396, -1416839988, -1103483252, 1052389004, -1103483252, -1103483252, 1065353216, -1103483252, 1044090914, -1162818823, -1103483252, -1416839988, -1166424545, 1044064338, -1103483252, -1416839988, 1049440636, -1111463718, -1235609300, -1093637749, 1058455711, -1103483252, -1103483250, 848972624, 1052389113, -1103472716, 958702290, 990013808, -1157455882, 1065353216, -1184696387, 962787261, -1103483252, -1103483252, -1288504488, 858979160, -1103483252, 1057727209, -1103477270, 951776135, -1103483252, -1416839988, 1057727209, -1103483251, 799198707, 1065353216, -1103483252, -1103483252, -1330688845, 816794803, -1183146888, 964336760, 1052389004, -1416839988, 1044000396, -1868328377, -1103483252, -1416839988, -1818962883, 1044000396, -1103483252, -1258026957, 1044022746, -1179755622, -1103483252, -1416821747, -1180849373, 1044020577, -1103483252, -1416839988, 1044000396, -1556267450, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044031480, -1175267368, -1103483252, -1261407310, -1103483252, -1173832630, 1044035426, -1416839988, -1627599725, -1103483252, 1044000396, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, -1103479293, 1044004355, -1321312984, -1416839988, -1392084868, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044133277, -1157512087, -1415904815, -1103483252, -1157536651, 1044132893, -1416839988, -1103483252, 1044055727, -1168628813, -1257866974, -1164097477, 1044080958, -1103483252, -1103483252, 1044000504, -1244025778, -1416839988, -1308784657, 1044000396, -1103483252, 1065353216, -1103483252, 1044000396, -1513223240, -1416839988, -1443694345, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044056342, -1168471584, -1416839988, -1103483252, -1189087920, 1044010633, -1211579584, -1103483252, 1044087299, -1163487040, -1416839988, -1166758063, 1044063035, -1103483252, 965537139, -1181946509, -1246912843, 900570805, 703736555, -1443747093, -1183743193, 963740455, 1065353216, -1263952095, 1044035432, -1173829724, -1103483252, -1416839988, -1175265170, 1044031484, -1103483252, -1416839988, 1044000396, -2078188789, -1103483252, -1416839988, -2005846931, 1044000396, -1103483252, -1103483252, 1044074949, -1164862337, -1416839988, -1165908946, 1044066772, -1103483252, -1103483252, 1044000396, -1531369661, -1416839988, -1599294534, 1044000396, -1103483252, -1258027103, 1044040337, -1172577290, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044000396, 0, -1103483252, -1416839988, -1103483252, 0, 1044000396, -1416821747, -1173055482, -1103483252, 1044038436, -1103483252, 1044000633, -1234332529, -1146889403, -1186176761, 1044349054, -1103483252, -1103483252, 1044012590, -1187084345, -1416839988, -1238420433, 1044000571, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044001116, -1221315657, -1283246431, -1103483252, -1171117794, 1044046009, -1283193683, -1103483252, 1044739686, -1137410719, -1416839988, -1139515844, 1044608111, -1103483252, -1103483252, 1044003208, -1204829201, -1146925620, -1176544024, 1044363432, -1103483252, 1065353216, -1103483252, 1044000481, -1247063573, -1416839988, -1308558949, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1353784249, -1065913784, -1103483252, -1298278099, 1082231448, -1166893263, -1103483252, 1044132807, -1165406652, -1398399119, -1168272552, 1044057119, -1103483252, -1176734614, 970749034, 967528232, -1179955416, -1249343934, 898139714, -1189281617, 958202031, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, -1189690414, 957793234, 846063501, -1301420147, 1063828015, -1103483252, -1103483252, -1103483252, -1103483252, 959290874, -1188192774, 973741937, -1173741711, 1060777612, -1103483252, -1103483252, -1323531519, 823952129, -1174084621, 973399027, -1103483252, -1103483252, 1060777612, -1214102462, 933381186, -1556299808, 591183840, -1200815871, 946667777, -1103483252, -1103483252, 0, 0, 1052389004, -1291371774, 856111874, -1182987271, 964496377, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, 328353268, -1819130380, 946667489, -1200816159, 141595410, -2005888238, -1197802529, 949681119, -1534506417, 612977231, -1221665183, 925818465, 1052389004, 937122730, -1210360918, 0, 0, 0, 0, -1239934895, 907548753, -1103483252, -1103483252, -1103483252, 1057727209, -1103483252, 802209880, -1103485389, -1207173495, 1085283848, -1103483252, 722622313, -1103483251, 846626608, -1416839988, -1416839988, 905994125, -1239781880, -1103483021, 912766372, 954183752, -1193231045, -1103471564, 959881826, -1190552070, 954272549, -1239641937, 906452166, -1103480035, 944312925, -1416839988, -1416839988, -1103492781, -1189809184, -1161175527, 986307593, -1103483253, -1065913784, -1166003173, 945590342, 1065353216, -1103479758, 945446711, -1103483252, -1416839988, 1075309154, -1103483257, -1281483635, -1103476928, 952476548, -1218853170, 928089673, -1416839988, -1416839988, -1103483252, -1416839988, -1103479293, 805636190, -1103483231, 883703842, -1103483252, -1416839988, -1416839988, -1416839988, -1103483252, -1416840177, -1214894333, 932318917, -1103484984, -1146834005, -1103480883, 940842127, -1103487103, -1146802399, -1103483235, 881272503, 1065353216, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103483252, -1103483252, -1103483252, 968153757, -1179329891, -1196443316, 951040332, -1103483252, 1060777612, 191506128, -1955977520, -1481862849, 665620799, -1228682415, 918801233, -1188398473, 959085175, -1103483252, -1103483252, 1052389004, 0, 0, 890643247, -1256840401, 951730480, -1195753168, -1183937866, 963545782, -1103483252, -1103483252, 693303474, -1454180174, 1050626690, -1096856958, 1052389004, -1103482945, 916040913, 1071289810, -1103491760, -1111775831, -1103483257, -1243143682, -1087044365, 790348910, -1103480791, 941217859, -1103478006, 950268365, -1192537452, 954946112, 1065353216, -1103483252, -1416839988, 940496387, -1206987256, -1103483252, -1416863964, -1103483252, -1416839988, 1070522257, -1103479852, 945064316, 877692018, -1087044362, -1103492407, -1190196732, 1065353216, 868543751, -1278939897, -1404663328, 742820320, 869407191, -1278076457, -1404660202, 742823446, 868835333, -1278648315, -1404807612, 742676036, 867962261, -1279521387, -1404656520, 742827128, 869211464, -1278272184, -1404660388, 742823260, 868329071, -1279154577, -1404623085, 742860563, 869201539, -1278282109, -1404660374, 742823274, 869216915, -1278266733, -1404657402, 742826246, 1065353216, -1416839988, 1044000396, -1680870018, -1103483252, -1416839988, -1631766710, 1044000396, -1103483252, -1416839988, 1044009553, -1190194069, -1103483252, -1280845202, -1181738849, 1044018845, -1103483252, -1103483252, 1044113763, -1159894129, -1414234099, -1159914818, 1044113601, -1103483252, -1103483252, 1044000396, -1572552438, -1416839988, -1641111818, 1044000396, -1103483252, -1103483252, 1044000396, -1610467424, -1416839988, -1669184958, 1044000396, -1103483252, -1103483252, 1044025499, -1178329567, -1416839988, -1184732988, 1044014886, -1103483252, 1044000396, 0, -1103483252, 0, 1071755232, -1077253617, -1103483252, 1044089771, -1162965132, -1103483252, -1163353941, 1044086733, -1416839913, -1103483252, 1044000396, -1750925261, -1103483252, -1686985275, 1044000396, -1416839988, -1103483252, 1065353216, -1103483252, 1044000396, -1416839988, 1044000396, -1103483252, -1103483252, 1052389004, -1103483252, -1416839988, -1103483252, 1044000496, -1245180522, -1065913784, -1184996871, 1082231893, -1103483252, 1052389004, -1103483252, -1103483252, 1044014306, -1185326941, -1103483252, -1103483252, -1238890911, 1044000564, -1416839988, -1103483252, 1044000396, -2147483647, -1416839988, -2147483147, 1044000396, -1416839988, -1103483252, 1065353216, -1103483252, 1044000910, -1224699803, -1125448600, -1183881047, 1045940979, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1708300623, -1416839988, -1103483252, -1765887542, 1044000396, -1416839171, -1103483252, 1044057492, -1168177009, -1296226300, -1166648854, 1044063463, -1103483252, -1103483252, 1044000546, -1240036050, -1173114061, -1181467364, 1044057181, -1103483252, -1103483252, 1044008643, -1191125278, -1416839988, -1245430777, 1044000494, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044041060, -1172383691, -1416839749, -1103483252, -1173307327, 1044037452, -1065913784, -1103483252, 1082232357, -1176289335, -1416839988, -1214941355, 1044001591, -1103483252, -1103483252, -1103483252, -1207620341, 939863307, 1052389004, -1103483252, -1103483252, 947016362, -1200467286, -1178570314, 968913334, 1052389004, 0, 0, -1220097516, 927386132, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, -1103481010, 940320411, -1103480519, 942329935, -1416839988, -1416839988, 1083816814, -1103485351, -1125431814, -1103481587, 936386447, -1103481775, 934847568, -1065913581, 944485613, 1065353216, -1103483252, -1077253617, -1103483252, -1416839988, 1087074187, -1103483252, -1416839988, 941082365, -1065913632, -1103483252, -1416839988, 939705092, -1207772503, -1103483831, -1172965871, 1065353216, -1616579275, 530904373, -1193466441, 954017207, -1103483252, -1103483252, 1052389004, -1103483252, -1103483252, -1188297610, 959186038, -1713869634, 433614014, 965642821, -1181840827, -1194679056, 952804592, 1052389004, -1103483252, -1103483252, -1103483252, -1103483252, 1060777612, 546261305, -1601222343, 967907670, -1179575978, -1103483252, -1103483252, 460414917, -1687068731, 959897630, -1187586018, 499, -2147483149, 960927468, -1186556180, 1052389004, -1416839988, 1044000396, -1955527681, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1382098153, 1044030485, -1175776537, -1103483252, -1416839987, -1103483252, -1179739628, 1044022745, -1416839988, -1895536330, -1103483252, 1044000396, -1103483252, 1044001288, -1218500854, -1234116533, -1177552844, 1044027257, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044113665, -1159906646, -1414508673, -1103483252, -1159934427, 1044113448, -1414525614, -1103483252, 1044085082, -1163565277, -1246169173, -1162425846, 1044094076, -1103483252, -1103483252, 1044000508, -1243502471, -1416839988, -1308389027, 1044000396, -1103483252, 1065353216, -1103483252, 1044004426, -1199841244, -1234159908, -1172213951, 1044041963, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044030642, -1175696274, -1416839988, -1103483252, -1238429260, 1044000571, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, 951700825, -1195782823, -1246495935, 900987713, 971327885, -1176155763, 0, 0, 1065353216, -1314070729, 1044462120, -1142852735, -1103483252, -1416839988, -1181167240, 1044019956, -1103483252, -1416839988, 1044000484, -1246714995, -1103483252, -1234120428, -1194043659, 1044007431, -1103483252, -1103483252, 1044085170, -1163553991, -1415753253, -1163615452, 1044084690, -1103483252, -1103483252, 1044000396, -1530696379, -1416839988, -1599140746, 1044000396, -1103483252, -1416839988, 1044009540, -1190206813, -1103483252, 1052389339, -1103483252, -1103483252, -1222130260, -1416839988, 1044000396, -1631111446, -1103483252, -1416839988, -1103483252, -1680149846, 1044000396, -1281158280, -1181743035, -1103483252, 1044018837, -1103483252, 1044046457, -1171002095, -1355359350, -1170725880, 1044047536, -1103483252, -1103483252, 1044000396, -1979167291, -1416839988, -1909069008, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, -1641926248, -1416839988, -1103483252, -1703575569, 1044000396, -1416839988, -1103483252, 1044033941, -1174206151, -1416839988, -1234337217, 1044000633, -1103483252, -1103483252, 1044000429, -1257989115, -1354357725, -1209069219, 1044002308, -1103483252, 1065353216, -1103483252, 1044000508, -1243569610, -1416839988, -1308429492, 1044000396, -1103483252, 1052389004, -1103483252, -1103483252, -1103483252, 1044000396, 0, -1416839988, -1103483252, 0, 1044000396, -1416839988, -1103483252, 1044000396, 0, -1416839988, 0, 1044000396, -1103483252, -1178479308, 969004340, 935529521, -1211954127, -1246549518, 900934130, 0, 0, 1065353216, -1222130260, -1103483252, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, 923524850, -1223958798, -1647615706, 499867942, 1060777612, 953317977, -1194165671, 250675443, -1896808205, -1147204443, 1000279205, -1103483252, -1103483252, -1631335648, 516148000, 1052389004, -1103483252, -1103483252, 967429273, -1180054375, -1180829381, 966654267, -1103483252, -1103483252, 1060777612, -1103483252, 695803022, -1451680626, -1177433330, 970050318, -1222130260, -1103483252, -1103483252, 1057727376, -1103483252, -1103483252, -1103483252, -1103483252, -1103483252, 238379747, -1909103901, 0, 0, 1063828015, -1582779429, 564704219, -1246814899, 900668749, -1575973942, 571509706, -1242873905, 904609743, -1103483252, -1103483252, -1103483252, 1057727209, -1103483252, -1416707932, 1070691433, -1103483252, 722945600, -1416839988, -1416839988, -1103483178, 898901971, -1103483252, -1416839988, -1208312334, 939171304, -1103483153, 902222364, 943243809, -1203861025, -1103473402, 957999647, -1416839988, -1416839988, -1159502019, 987981585, -1103483046, 911083953, -1416839988, -1416839988, -1103483252, -1416839988, -1190869900, 956613748, -1103483252, -1416839988, -1416839988, -1416839988, 1065353216, -1103483252, -1416839992, -1103474590, 956782682, 1075267071, -1103483258, -1281035152, 941588119, -1205874043, -1103483252, -1416839994, -1103479716, 945619596, -1416839988, -1416839988, -1103487246, -1199288178, -1103483230, 884119604, -1103491201, -1191189131, 931508748, -1214002129, -1103483252, -1416840187, 941589190, -1205873584, -1103483772, -1224614051, -1103483252, -1416839988, -1103483571, -1231060292, -1103483230, 884066643, 1065353216, -1103483252, -1103483252, 515503988, -1631979660, -1196213294, 951270354, 951068643, -1196415005, -1232531452, 914952196, -1534006351, 613477297, 953326187, -1194157461, 1052389004};
localparam integer A_BRAMInd[0:5851] = '{0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 3, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 3, 1, 2, 3, 0, 3, 0, 3, 0, 1, 2, 3, 3, 0, 3, 0, 1, 2, 2, 1, 2, 3, 3, 0, 1, 1, 2, 2, 0, 2, 3, 1, 2, 1, 3, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 1, 3, 0, 3, 0, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 1, 2, 1, 0, 0, 1, 2, 3, 1, 2, 3, 2, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 0, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 1, 2, 2, 1, 2, 3, 0, 1, 2, 3, 0, 2, 2, 3, 2, 2, 3, 1, 3, 3, 0, 3, 0, 0, 1, 2, 1, 1, 2, 1, 1, 2, 3, 2, 2, 3, 2, 2, 3, 0, 3, 0, 0, 1, 0, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 2, 3, 1, 2, 3, 0, 1, 3, 0, 1, 2, 1, 1, 2, 0, 1, 0, 1, 2, 3, 1, 1, 2, 3, 2, 3, 1, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 3, 1, 3, 1, 2, 3, 0, 1, 2, 3, 0, 0, 2, 3, 3, 1, 2, 3, 1, 2, 1, 2, 3, 0, 1, 0, 1, 2, 3, 0, 2, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 3, 0, 1, 2, 0, 1, 2, 3, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 1, 3, 0, 1, 2, 3, 0, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 0, 2, 3, 0, 1, 3, 3, 0, 2, 3, 0, 1, 3, 0, 3, 0, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 0, 1, 0, 2, 3, 2, 0, 1, 2, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 0, 1, 2, 1, 0, 1, 2, 0, 1, 2, 0, 2, 3, 0, 1, 2, 3, 0, 1, 0, 2, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 0, 1, 2, 1, 3, 1, 2, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 2, 0, 1, 0, 2, 3, 0, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 3, 0, 3, 1, 2, 1, 3, 0, 1, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 2, 3, 3, 1, 2, 1, 3, 0, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 2, 0, 1, 3, 1, 3, 0, 3, 1, 2, 0, 2, 3, 0, 1, 1, 0, 1, 3, 1, 3, 0, 3, 1, 0, 1, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 2, 0, 1, 0, 2, 3, 0, 1, 2, 3, 0, 2, 1, 2, 0, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 1, 0, 1, 2, 3, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 3, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 0, 2, 3, 0, 1, 3, 0, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 3, 1, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 3, 0, 3, 1, 3, 0, 1, 2, 2, 2, 0, 2, 3, 0, 1, 0, 1, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 2, 3, 0, 1, 3, 2, 3, 0, 3, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 0, 0, 1, 2, 3, 2, 3, 0, 1, 0, 1, 2, 0, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 2, 3, 3, 2, 3, 2, 3, 0, 1, 1, 2, 1, 2, 1, 3, 0, 2, 3, 0, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 2, 0, 1, 2, 3, 1, 3, 0, 1, 2, 3, 0, 3, 0, 1, 2, 3, 0, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 3, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 0, 2, 3, 0, 1, 2, 3, 3, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 2, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 2, 3, 2, 0, 2, 3, 0, 1, 0, 1, 3, 1, 2, 3, 0, 3, 0, 1, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 1, 3, 2, 3, 0, 1, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 0, 0, 1, 2, 3, 2, 3, 0, 1, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 0, 1, 3, 1, 3, 0, 1, 2, 3, 0, 2, 2, 0, 1, 0, 1, 3, 0, 3, 0, 3, 0, 3, 0, 1, 3, 0, 1, 2, 0, 1, 2, 0, 2, 3, 1, 2, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 2, 3, 0, 1, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 0, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 3, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 0, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 1, 3, 0, 1, 2, 3, 0, 0, 3, 0, 1, 2, 3, 0, 1, 2, 1, 0, 1, 2, 0, 1, 3, 0, 3, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 0, 1, 3, 3, 2, 3, 1, 0, 1, 2, 0, 3, 0, 2, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 0, 1, 3, 2, 3, 0, 2, 3, 2, 3, 1, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 3, 0, 1, 2, 3, 1, 0, 1, 2, 0, 3, 0, 1, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 1, 0, 1, 2, 0, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 1, 2, 0, 0, 3, 0, 2, 1, 2, 3, 1, 0, 1, 3, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 1, 2, 0, 3, 0, 1, 3, 0, 3, 0, 2, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 2, 3, 2, 0, 2, 3, 0, 1, 1, 2, 0, 2, 3, 0, 1, 0, 1, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 2, 3, 0, 1, 3, 2, 3, 0, 3, 3, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 1, 1, 2, 3, 0, 3, 0, 1, 2, 1, 2, 3, 1, 1, 2, 3, 0, 2, 3, 0, 1, 2, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 3, 0, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 1, 3, 0, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 0, 1, 1, 2, 1, 2, 3, 1, 2, 0, 1, 2, 3, 1, 2, 3, 1, 3, 0, 2, 3, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 2, 3, 0, 1, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 1, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 2, 0, 1, 2, 3, 0, 1, 1, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 3, 2, 3, 0, 1, 2, 3, 0, 1, 3, 1, 2, 1, 3, 0, 1, 3, 0, 3, 3, 0, 1, 2, 2, 1, 2, 1, 2, 3, 0, 1, 2, 3, 1, 0, 1, 2, 3, 0, 1, 2, 3, 2, 2, 3, 0, 1, 3, 0, 1, 2, 0, 0, 3, 0, 1, 2, 3, 0, 3, 2, 2, 3, 0, 1, 3, 1, 2, 3, 2, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 3, 1, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 1, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 3, 0, 1, 2, 3, 0, 1, 2, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 1, 2, 1, 0, 2, 3, 0, 1, 2, 3, 0, 2, 1, 2, 1, 2, 0, 1, 1, 2, 1, 2, 1, 3, 0, 2, 3, 0, 1, 3, 1, 3, 0, 1, 2, 0, 1, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 1, 2, 3, 0, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 1, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 2, 0, 1, 2, 3, 0, 1, 1, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 1, 2, 3, 1, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 0, 1, 2, 0, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 2, 0, 1, 2, 0, 1, 2, 3, 0, 1, 3, 0, 1, 1, 0, 1, 0, 2, 3, 1, 2, 3, 3, 3, 1, 3, 0, 1, 2, 1, 2, 1, 1, 2, 3, 0, 1, 2, 3, 0, 2, 2, 3, 0, 1, 3, 2, 3, 0, 0, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 2, 2, 3, 0, 1, 3, 0, 1, 2, 1, 3, 0, 2, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 1, 2, 0, 1, 2, 1, 3, 0, 2, 3, 2, 2, 1, 2, 1, 2, 0, 1, 1, 2, 1, 2, 2, 0, 1, 3, 0, 1, 2, 1, 2, 3, 1, 3, 0, 2, 3, 3, 1, 2, 3, 0, 1, 2, 3, 0, 2, 0, 1, 3, 0, 1, 2, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 0, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 1, 3, 0, 1, 2, 3, 0, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 3, 1, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 3, 0, 3, 1, 3, 0, 1, 2, 3, 2, 0, 2, 3, 0, 1, 0, 1, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 0, 3, 0, 1, 3, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 3, 3, 0, 1, 2, 1, 2, 3, 0, 3, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 3, 0, 2, 1, 3, 0, 1, 2, 3, 0, 2, 2, 1, 2, 1, 2, 0, 1, 0, 1, 0, 1, 1, 3, 0, 2, 3, 0, 1, 3, 0, 1, 3, 1, 2, 0, 1, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 1, 2, 3, 0, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 2, 3, 0, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 1, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 3, 0, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 1, 3, 0, 1, 2, 3, 0, 3, 1, 2, 3, 0, 0, 1, 0, 1, 2, 3, 3, 1, 2, 3, 0, 1, 3, 0, 1, 2, 2, 0, 2, 3, 1, 2, 3, 0, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 1, 2, 3, 1, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 0, 1, 2, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 2, 3, 0, 1, 3, 0, 3, 1, 3, 0, 1, 2, 1, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 3, 0, 2, 1, 2, 3, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 2, 3, 2, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 1, 2, 3, 0, 3, 0, 3, 0, 1, 0, 1, 2, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 2, 0, 1, 2, 3, 2, 3, 0, 2, 3, 0, 1, 2, 3, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 3, 1, 2, 3, 0, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 0};
localparam integer A_BRAMAddr[0:5851] = '{0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 7, 7, 7, 8, 8, 8, 9, 9, 9, 9, 10, 10, 10, 10, 11, 11, 11, 11, 12, 12, 12, 12, 13, 13, 13, 13, 14, 14, 14, 14, 15, 15, 15, 15, 16, 16, 16, 16, 17, 17, 18, 18, 18, 18, 19, 19, 19, 19, 20, 20, 20, 20, 21, 21, 21, 21, 22, 22, 22, 22, 23, 23, 23, 23, 24, 24, 24, 24, 25, 25, 25, 25, 26, 26, 26, 26, 27, 27, 27, 27, 28, 28, 28, 29, 29, 29, 30, 30, 30, 30, 31, 31, 32, 32, 32, 32, 33, 33, 33, 33, 34, 34, 34, 34, 35, 35, 35, 35, 36, 36, 36, 36, 37, 37, 37, 37, 38, 38, 38, 38, 39, 39, 39, 39, 40, 40, 40, 40, 41, 41, 41, 41, 42, 42, 42, 42, 43, 43, 43, 44, 44, 44, 45, 45, 45, 45, 46, 46, 46, 46, 47, 47, 47, 47, 48, 48, 48, 48, 49, 49, 49, 49, 50, 50, 50, 51, 51, 51, 52, 52, 52, 52, 53, 53, 53, 53, 54, 54, 54, 54, 55, 55, 55, 55, 56, 56, 56, 56, 57, 57, 57, 57, 58, 58, 58, 58, 59, 59, 59, 60, 60, 60, 61, 61, 61, 61, 62, 62, 62, 63, 63, 64, 64, 64, 65, 65, 65, 66, 66, 66, 66, 67, 67, 68, 68, 68, 69, 69, 69, 69, 70, 70, 70, 70, 71, 71, 71, 71, 72, 72, 72, 73, 74, 74, 74, 74, 75, 75, 75, 76, 76, 76, 76, 77, 77, 77, 77, 78, 79, 79, 79, 80, 80, 81, 81, 83, 83, 83, 83, 84, 85, 85, 86, 86, 86, 87, 88, 88, 88, 89, 90, 90, 91, 91, 92, 93, 93, 93, 94, 94, 95, 95, 96, 96, 97, 97, 97, 97, 98, 98, 98, 98, 99, 99, 100, 100, 101, 101, 102, 102, 103, 103, 103, 103, 104, 104, 104, 104, 105, 105, 105, 105, 106, 106, 106, 106, 107, 107, 107, 107, 108, 108, 108, 108, 109, 109, 109, 109, 110, 111, 111, 112, 113, 114, 114, 114, 114, 115, 115, 115, 116, 117, 117, 117, 118, 118, 118, 118, 119, 120, 120, 121, 122, 122, 122, 123, 123, 123, 124, 124, 124, 124, 125, 125, 125, 125, 126, 126, 126, 126, 127, 127, 127, 127, 128, 128, 128, 128, 129, 129, 129, 129, 130, 130, 130, 131, 131, 131, 132, 132, 132, 132, 133, 133, 133, 133, 134, 134, 134, 135, 135, 135, 136, 136, 136, 136, 137, 137, 137, 138, 138, 138, 138, 139, 139, 139, 139, 140, 140, 140, 140, 141, 141, 142, 142, 142, 142, 143, 143, 143, 144, 144, 144, 144, 145, 145, 146, 147, 147, 147, 148, 148, 148, 148, 149, 149, 150, 150, 151, 152, 152, 153, 153, 154, 155, 155, 156, 157, 157, 157, 158, 159, 159, 160, 161, 161, 161, 162, 163, 163, 164, 165, 165, 166, 166, 167, 168, 168, 169, 170, 170, 170, 171, 171, 171, 171, 172, 172, 172, 172, 173, 173, 173, 174, 174, 174, 175, 175, 175, 175, 176, 176, 176, 176, 177, 177, 177, 178, 179, 179, 180, 180, 181, 181, 181, 181, 182, 182, 182, 182, 183, 183, 183, 184, 185, 185, 186, 187, 187, 188, 188, 188, 189, 189, 189, 190, 191, 191, 192, 192, 193, 193, 193, 193, 194, 195, 195, 195, 196, 196, 197, 198, 198, 198, 198, 199, 199, 200, 200, 200, 200, 202, 202, 202, 202, 203, 204, 205, 205, 205, 206, 207, 208, 208, 208, 209, 209, 209, 209, 210, 212, 212, 212, 213, 214, 214, 214, 215, 215, 217, 217, 217, 218, 218, 219, 219, 219, 219, 220, 220, 221, 221, 221, 221, 223, 223, 224, 224, 224, 224, 225, 225, 225, 225, 226, 226, 226, 226, 227, 227, 227, 228, 228, 229, 229, 229, 230, 230, 230, 230, 231, 231, 232, 232, 232, 233, 233, 233, 233, 234, 236, 236, 236, 237, 237, 237, 237, 238, 238, 238, 238, 239, 239, 240, 240, 240, 241, 241, 241, 241, 242, 242, 243, 243, 243, 244, 244, 244, 244, 245, 245, 245, 245, 246, 246, 246, 248, 248, 249, 249, 249, 249, 250, 250, 250, 250, 251, 251, 251, 251, 252, 252, 252, 252, 253, 253, 253, 253, 254, 254, 254, 254, 255, 255, 255, 255, 256, 256, 256, 256, 257, 257, 257, 257, 258, 258, 258, 259, 259, 259, 260, 260, 260, 260, 261, 261, 261, 261, 262, 262, 262, 262, 263, 263, 263, 263, 264, 264, 264, 264, 265, 265, 265, 265, 266, 266, 266, 267, 267, 267, 267, 268, 268, 269, 269, 269, 269, 270, 270, 270, 271, 271, 271, 272, 272, 272, 273, 274, 274, 274, 275, 275, 275, 276, 277, 278, 278, 278, 280, 280, 280, 281, 281, 281, 281, 282, 282, 282, 282, 283, 283, 283, 283, 284, 284, 284, 284, 285, 285, 285, 285, 286, 286, 286, 286, 287, 287, 287, 288, 288, 288, 289, 289, 289, 289, 290, 290, 290, 290, 291, 291, 291, 291, 292, 292, 292, 292, 293, 293, 293, 293, 294, 294, 294, 294, 295, 295, 295, 295, 296, 296, 296, 297, 297, 297, 298, 298, 298, 298, 299, 299, 299, 299, 300, 300, 300, 300, 301, 301, 301, 301, 302, 302, 302, 302, 303, 303, 303, 303, 304, 304, 304, 304, 305, 305, 306, 306, 306, 306, 307, 307, 307, 308, 308, 309, 309, 309, 310, 311, 311, 311, 312, 312, 312, 312, 313, 313, 313, 314, 314, 314, 314, 315, 315, 315, 315, 316, 316, 316, 316, 317, 317, 317, 317, 318, 318, 318, 318, 319, 319, 319, 319, 320, 320, 320, 320, 321, 321, 321, 321, 322, 323, 323, 323, 323, 324, 324, 324, 324, 325, 325, 325, 326, 326, 326, 327, 327, 327, 327, 328, 328, 328, 328, 329, 329, 329, 329, 330, 330, 330, 330, 331, 331, 331, 331, 332, 332, 332, 332, 333, 333, 333, 333, 334, 334, 334, 334, 335, 335, 335, 335, 336, 336, 336, 336, 337, 337, 337, 338, 338, 338, 339, 339, 339, 339, 340, 340, 340, 340, 341, 341, 341, 341, 342, 342, 342, 342, 343, 343, 343, 343, 344, 344, 344, 344, 345, 345, 345, 345, 346, 346, 346, 347, 347, 347, 348, 348, 348, 348, 349, 349, 349, 349, 350, 350, 350, 350, 351, 351, 351, 351, 352, 352, 352, 352, 353, 353, 353, 353, 354, 354, 354, 355, 355, 355, 356, 356, 356, 356, 357, 357, 357, 358, 358, 359, 359, 359, 360, 361, 361, 361, 362, 362, 362, 363, 363, 363, 364, 364, 364, 364, 365, 365, 366, 366, 367, 367, 367, 368, 368, 368, 369, 369, 369, 369, 370, 370, 370, 370, 371, 371, 371, 371, 372, 372, 372, 372, 373, 373, 374, 374, 375, 375, 375, 376, 376, 377, 377, 377, 378, 378, 379, 379, 380, 380, 380, 381, 381, 381, 381, 382, 382, 382, 382, 383, 383, 383, 383, 384, 384, 384, 384, 385, 385, 385, 385, 386, 386, 386, 386, 387, 387, 387, 387, 388, 388, 388, 388, 389, 389, 389, 389, 390, 390, 390, 391, 391, 391, 392, 392, 392, 392, 393, 393, 393, 393, 394, 394, 394, 394, 395, 395, 395, 395, 396, 396, 396, 396, 397, 397, 397, 397, 398, 398, 398, 398, 399, 399, 399, 400, 400, 400, 401, 401, 401, 401, 402, 402, 402, 402, 403, 403, 403, 403, 404, 404, 404, 404, 405, 405, 405, 405, 406, 406, 406, 406, 407, 407, 407, 407, 408, 408, 408, 409, 409, 409, 410, 410, 410, 410, 411, 411, 411, 412, 413, 413, 414, 414, 414, 415, 415, 415, 416, 416, 416, 417, 417, 417, 417, 418, 418, 418, 418, 419, 419, 420, 420, 420, 420, 421, 421, 421, 421, 422, 422, 422, 422, 423, 423, 423, 423, 424, 424, 424, 424, 425, 425, 425, 425, 426, 426, 426, 426, 427, 427, 427, 427, 428, 428, 429, 429, 429, 429, 430, 430, 430, 430, 431, 431, 431, 431, 432, 432, 432, 432, 433, 433, 433, 433, 434, 434, 434, 434, 435, 435, 435, 435, 436, 436, 436, 437, 437, 437, 438, 438, 438, 438, 439, 439, 439, 440, 440, 441, 441, 442, 442, 443, 443, 443, 444, 444, 444, 445, 445, 445, 445, 446, 446, 446, 446, 447, 447, 447, 447, 448, 448, 448, 448, 449, 449, 449, 449, 450, 450, 450, 450, 451, 451, 451, 451, 452, 452, 452, 452, 453, 453, 454, 454, 454, 455, 455, 455, 455, 456, 456, 456, 456, 457, 457, 458, 458, 458, 458, 459, 459, 459, 460, 460, 460, 460, 461, 461, 461, 461, 462, 463, 463, 463, 464, 464, 465, 466, 466, 467, 467, 468, 468, 469, 469, 469, 469, 470, 470, 470, 470, 471, 471, 471, 471, 472, 472, 472, 472, 473, 473, 473, 474, 474, 474, 475, 475, 475, 475, 476, 476, 476, 477, 478, 478, 478, 479, 479, 480, 480, 481, 481, 482, 482, 482, 483, 483, 484, 485, 485, 485, 486, 486, 487, 487, 488, 489, 489, 489, 490, 490, 491, 491, 491, 491, 492, 492, 492, 492, 493, 493, 493, 493, 494, 494, 494, 494, 495, 495, 495, 495, 496, 496, 496, 496, 497, 497, 497, 498, 498, 498, 499, 499, 499, 499, 500, 500, 500, 501, 502, 502, 503, 503, 503, 504, 504, 504, 504, 505, 505, 506, 506, 507, 507, 508, 508, 508, 509, 509, 509, 509, 510, 510, 510, 510, 511, 511, 511, 511, 512, 512, 512, 512, 513, 513, 513, 513, 514, 514, 514, 514, 515, 515, 515, 516, 517, 517, 517, 517, 518, 518, 518, 518, 519, 519, 519, 520, 520, 520, 521, 521, 521, 521, 522, 522, 522, 522, 523, 523, 523, 523, 524, 524, 524, 524, 525, 525, 525, 525, 526, 526, 526, 526, 527, 527, 527, 527, 528, 528, 528, 528, 529, 529, 529, 529, 530, 530, 530, 530, 531, 531, 531, 532, 532, 532, 533, 533, 533, 533, 534, 534, 534, 534, 535, 535, 535, 535, 536, 536, 536, 536, 537, 537, 537, 537, 538, 538, 538, 538, 539, 539, 539, 539, 540, 540, 541, 541, 541, 541, 542, 542, 542, 542, 543, 543, 543, 543, 544, 544, 544, 544, 545, 545, 545, 545, 546, 546, 546, 546, 547, 547, 547, 547, 548, 548, 548, 548, 549, 549, 550, 550, 550, 550, 551, 551, 551, 551, 552, 552, 553, 553, 554, 555, 555, 555, 555, 556, 556, 556, 557, 557, 558, 558, 558, 558, 559, 559, 559, 559, 560, 560, 560, 560, 561, 561, 561, 561, 562, 562, 562, 562, 563, 563, 563, 563, 564, 564, 564, 564, 565, 565, 565, 565, 566, 567, 567, 567, 567, 568, 568, 568, 568, 569, 569, 569, 570, 570, 570, 571, 571, 571, 571, 572, 572, 572, 572, 573, 573, 573, 573, 574, 574, 574, 574, 575, 575, 575, 575, 576, 576, 576, 576, 577, 577, 577, 577, 578, 578, 578, 578, 579, 579, 579, 579, 580, 580, 580, 580, 581, 581, 581, 581, 582, 582, 582, 582, 583, 583, 583, 583, 584, 584, 584, 584, 585, 585, 585, 585, 586, 586, 586, 586, 587, 587, 587, 587, 588, 588, 588, 588, 589, 589, 589, 589, 590, 590, 590, 590, 591, 591, 591, 591, 592, 592, 592, 592, 593, 593, 593, 594, 594, 594, 595, 595, 595, 595, 596, 596, 596, 596, 597, 597, 597, 598, 598, 598, 599, 599, 599, 600, 600, 601, 601, 601, 601, 602, 602, 602, 603, 603, 603, 604, 604, 604, 605, 606, 606, 606, 607, 607, 607, 607, 608, 608, 608, 609, 609, 609, 609, 610, 610, 610, 611, 611, 611, 611, 612, 612, 612, 612, 613, 613, 613, 613, 614, 614, 614, 614, 615, 616, 616, 616, 617, 617, 618, 618, 618, 618, 619, 619, 619, 619, 620, 620, 620, 620, 621, 621, 621, 621, 622, 622, 622, 622, 623, 623, 623, 624, 624, 624, 625, 625, 625, 625, 626, 626, 626, 626, 627, 627, 627, 627, 628, 628, 628, 628, 629, 629, 629, 629, 630, 630, 630, 630, 631, 631, 631, 631, 632, 632, 632, 633, 633, 633, 634, 634, 634, 634, 635, 635, 635, 635, 636, 636, 636, 636, 637, 637, 638, 638, 638, 638, 639, 639, 639, 640, 640, 640, 640, 641, 641, 641, 642, 642, 642, 642, 643, 643, 643, 643, 644, 644, 644, 644, 645, 645, 645, 645, 646, 646, 646, 646, 647, 647, 647, 647, 648, 648, 648, 648, 649, 649, 650, 650, 650, 651, 652, 652, 652, 652, 653, 653, 653, 653, 654, 654, 654, 654, 655, 655, 655, 655, 656, 656, 656, 656, 657, 657, 657, 657, 658, 658, 659, 659, 659, 659, 660, 660, 660, 660, 661, 661, 661, 661, 662, 662, 662, 662, 663, 663, 663, 663, 664, 664, 664, 664, 665, 665, 665, 665, 666, 666, 666, 667, 667, 667, 668, 668, 668, 668, 669, 669, 669, 669, 670, 670, 670, 670, 671, 671, 672, 672, 673, 673, 673, 674, 674, 674, 674, 675, 675, 675, 675, 676, 677, 677, 678, 678, 679, 679, 680, 680, 680, 681, 682, 683, 683, 683, 684, 684, 685, 685, 686, 687, 688, 688, 688, 688, 689, 689, 689, 689, 690, 691, 692, 692, 693, 693, 693, 694, 694, 695, 695, 696, 697, 697, 697, 697, 698, 698, 698, 699, 699, 699, 699, 700, 700, 702, 703, 703, 703, 703, 704, 704, 705, 705, 706, 706, 706, 707, 708, 708, 708, 708, 709, 709, 709, 709, 710, 710, 710, 711, 711, 711, 712, 712, 712, 712, 713, 713, 713, 713, 714, 714, 714, 714, 715, 715, 715, 716, 716, 716, 716, 717, 717, 719, 720, 720, 721, 721, 721, 721, 722, 722, 722, 723, 723, 723, 723, 724, 724, 724, 724, 725, 725, 725, 725, 726, 726, 726, 726, 727, 727, 727, 727, 728, 728, 728, 728, 729, 729, 731, 732, 732, 733, 733, 734, 735, 735, 736, 736, 737, 737, 738, 738, 739, 739, 740, 740, 741, 741, 741, 742, 742, 744, 744, 744, 745, 745, 745, 745, 746, 746, 747, 747, 747, 748, 748, 748, 748, 750, 750, 751, 751, 751, 751, 752, 752, 753, 753, 753, 753, 754, 754, 755, 755, 755, 756, 756, 756, 756, 757, 757, 757, 757, 758, 758, 759, 759, 761, 761, 762, 762, 762, 762, 763, 763, 763, 763, 764, 764, 764, 764, 765, 765, 765, 765, 766, 766, 766, 766, 767, 767, 767, 767, 768, 768, 768, 768, 769, 769, 769, 769, 770, 770, 770, 770, 771, 771, 771, 771, 772, 772, 772, 772, 773, 773, 773, 773, 774, 774, 774, 774, 775, 775, 775, 776, 776, 776, 777, 777, 777, 777, 778, 778, 778, 778, 779, 779, 779, 780, 780, 780, 781, 781, 781, 782, 782, 783, 783, 783, 783, 784, 784, 784, 785, 785, 785, 786, 786, 786, 786, 787, 788, 788, 788, 789, 789, 789, 789, 790, 790, 790, 791, 791, 791, 791, 792, 792, 792, 793, 793, 793, 793, 794, 794, 794, 794, 795, 795, 795, 795, 796, 796, 796, 797, 797, 798, 798, 799, 799, 799, 800, 800, 800, 800, 801, 801, 801, 801, 802, 802, 802, 802, 803, 803, 803, 803, 804, 804, 804, 804, 805, 805, 805, 806, 806, 806, 807, 807, 807, 807, 808, 808, 808, 808, 809, 809, 809, 809, 810, 810, 810, 810, 811, 811, 811, 811, 812, 812, 812, 812, 813, 813, 813, 813, 814, 814, 815, 815, 815, 815, 816, 816, 816, 816, 817, 817, 817, 817, 818, 818, 818, 819, 819, 819, 820, 820, 820, 820, 821, 821, 821, 822, 822, 822, 822, 823, 823, 823, 824, 824, 824, 824, 825, 825, 825, 825, 826, 826, 826, 826, 827, 827, 827, 827, 828, 828, 828, 828, 829, 829, 829, 829, 830, 830, 830, 830, 831, 832, 832, 832, 833, 833, 834, 834, 834, 834, 835, 835, 835, 835, 836, 836, 836, 836, 837, 837, 837, 837, 838, 838, 838, 838, 839, 839, 839, 840, 840, 840, 841, 841, 841, 841, 842, 842, 842, 842, 843, 843, 843, 843, 844, 844, 844, 844, 845, 845, 845, 845, 846, 846, 846, 846, 847, 847, 847, 847, 848, 848, 848, 849, 849, 849, 850, 850, 850, 850, 851, 851, 851, 851, 852, 852, 852, 852, 853, 853, 854, 854, 855, 855, 855, 856, 856, 856, 856, 857, 857, 857, 857, 858, 859, 859, 860, 861, 861, 861, 862, 862, 864, 864, 864, 865, 865, 865, 866, 866, 867, 868, 869, 869, 869, 869, 870, 870, 870, 870, 871, 871, 872, 873, 873, 874, 874, 874, 875, 875, 876, 876, 877, 877, 877, 877, 878, 878, 878, 879, 879, 879, 879, 880, 880, 880, 882, 883, 883, 883, 883, 884, 884, 885, 885, 886, 886, 886, 886, 888, 888, 889, 889, 889, 889, 890, 890, 890, 891, 891, 891, 891, 892, 892, 892, 893, 893, 893, 893, 894, 894, 894, 894, 895, 895, 895, 896, 896, 896, 896, 897, 897, 897, 897, 900, 901, 901, 901, 901, 902, 902, 902, 902, 903, 903, 903, 904, 904, 904, 904, 905, 905, 905, 905, 906, 906, 906, 906, 907, 907, 907, 907, 908, 908, 908, 908, 909, 909, 909, 909, 912, 913, 913, 914, 914, 914, 915, 915, 916, 916, 916, 916, 917, 917, 918, 919, 919, 920, 920, 920, 921, 921, 922, 922, 923, 923, 925, 925, 925, 926, 926, 926, 927, 927, 927, 928, 928, 928, 929, 929, 930, 931, 931, 931, 931, 932, 932, 932, 932, 933, 933, 934, 934, 934, 935, 935, 936, 937, 937, 937, 938, 938, 938, 938, 939, 939, 939, 939, 940, 940, 941, 941, 943, 943, 943, 944, 944, 944, 944, 945, 945, 946, 946, 946, 947, 947, 948, 948, 948, 949, 949, 949, 949, 950, 950, 950, 950, 951, 951, 951, 951, 952, 952, 952, 952, 953, 953, 953, 953, 954, 954, 954, 954, 955, 955, 955, 955, 956, 956, 956, 956, 957, 957, 957, 957, 958, 958, 958, 959, 959, 959, 960, 960, 960, 960, 961, 961, 961, 961, 962, 962, 962, 962, 963, 963, 964, 964, 964, 965, 965, 965, 966, 966, 966, 967, 967, 967, 967, 968, 968, 969, 969, 969, 969, 970, 971, 971, 972, 972, 972, 972, 973, 973, 973, 974, 975, 975, 975, 976, 976, 976, 977, 977, 978, 978, 979, 979, 979, 980, 980, 980, 980, 981, 981, 981, 981, 982, 982, 983, 984, 984, 984, 985, 986, 986, 987, 988, 988, 988, 989, 989, 990, 990, 991, 991, 991, 992, 992, 992, 993, 993, 993, 993, 994, 994, 994, 995, 995, 995, 996, 996, 996, 996, 997, 997, 998, 998, 998, 999, 999, 1000, 1000, 1000, 1001, 1001, 1002, 1003, 1003, 1003, 1004, 1004, 1004, 1004, 1005, 1005, 1005, 1005, 1006, 1006, 1006, 1007, 1007, 1007, 1008, 1008, 1008, 1008, 1009, 1009, 1009, 1009, 1010, 1010, 1010, 1010, 1011, 1012, 1012, 1012, 1012, 1013, 1013, 1013, 1013, 1014, 1015, 1015, 1015, 1016, 1016, 1017, 1017, 1018, 1018, 1018, 1018, 1019, 1019, 1019, 1019, 1020, 1020, 1021, 1022, 1022, 1022, 1023, 1023, 1024, 1024, 1024, 1025, 1025, 1025, 1025, 1026, 1026, 1026, 1026, 1027, 1027, 1027, 1028, 1029, 1029, 1030, 1031, 1031, 1032, 1032, 1033, 1033, 1033, 1034, 1035, 1035, 1035, 1036, 1036, 1037, 1037, 1037, 1038, 1038, 1038, 1038, 1039, 1039, 1039, 1039, 1040, 1040, 1041, 1041, 1041, 1041, 1042, 1042, 1042, 1043, 1043, 1044, 1044, 1045, 1045, 1045, 1046, 1046, 1047, 1047, 1048, 1048, 1048, 1049, 1049, 1049, 1050, 1050, 1050, 1050, 1051, 1051, 1051, 1052, 1052, 1052, 1053, 1053, 1053, 1053, 1054, 1054, 1054, 1054, 1055, 1055, 1055, 1055, 1056, 1056, 1057, 1058, 1058, 1058, 1058, 1059, 1059, 1060, 1060, 1060, 1060, 1061, 1061, 1061, 1062, 1063, 1063, 1064, 1065, 1065, 1065, 1066, 1066, 1067, 1068, 1069, 1069, 1069, 1070, 1070, 1071, 1071, 1072, 1073, 1074, 1074, 1074, 1074, 1075, 1075, 1075, 1075, 1076, 1077, 1078, 1078, 1079, 1079, 1079, 1080, 1080, 1081, 1081, 1082, 1083, 1083, 1083, 1084, 1084, 1084, 1085, 1085, 1085, 1085, 1086, 1086, 1086, 1088, 1089, 1089, 1089, 1090, 1090, 1091, 1091, 1091, 1092, 1092, 1092, 1093, 1094, 1094, 1094, 1095, 1095, 1095, 1096, 1096, 1096, 1097, 1097, 1097, 1097, 1098, 1098, 1098, 1099, 1099, 1099, 1099, 1100, 1100, 1100, 1100, 1101, 1101, 1101, 1102, 1102, 1102, 1102, 1103, 1103, 1103, 1103, 1106, 1107, 1107, 1107, 1107, 1108, 1108, 1108, 1109, 1109, 1110, 1110, 1110, 1110, 1111, 1111, 1111, 1111, 1112, 1112, 1112, 1112, 1113, 1113, 1113, 1113, 1114, 1114, 1114, 1114, 1115, 1115, 1115, 1115, 1116, 1116, 1118, 1119, 1119, 1120, 1120, 1121, 1122, 1123, 1123, 1123, 1124, 1124, 1124, 1124, 1125, 1126, 1126, 1127, 1127, 1128, 1128, 1129, 1129, 1130, 1130, 1131, 1132, 1132, 1133, 1133, 1133, 1133, 1134, 1134, 1134, 1135, 1135, 1136, 1136, 1136, 1137, 1138, 1138, 1138, 1139, 1139, 1139, 1139, 1140, 1140, 1141, 1141, 1141, 1141, 1142, 1142, 1143, 1143, 1144, 1144, 1144, 1144, 1145, 1145, 1145, 1145, 1146, 1146, 1146, 1146, 1147, 1147, 1148, 1149, 1149, 1149, 1150, 1150, 1150, 1150, 1151, 1151, 1151, 1151, 1152, 1152, 1152, 1152, 1153, 1153, 1153, 1153, 1154, 1154, 1154, 1154, 1155, 1155, 1155, 1155, 1156, 1156, 1156, 1156, 1157, 1157, 1157, 1157, 1158, 1159, 1159, 1159, 1159, 1160, 1160, 1160, 1160, 1161, 1161, 1161, 1162, 1162, 1162, 1163, 1163, 1163, 1164, 1164, 1164, 1164, 1165, 1165, 1165, 1165, 1166, 1166, 1166, 1166, 1167, 1167, 1167, 1167, 1168, 1168, 1168, 1168, 1169, 1169, 1169, 1169, 1170, 1170, 1170, 1170, 1171, 1171, 1171, 1171, 1172, 1172, 1172, 1172, 1173, 1173, 1173, 1173, 1174, 1174, 1174, 1174, 1175, 1175, 1175, 1175, 1176, 1176, 1176, 1176, 1177, 1177, 1177, 1177, 1178, 1178, 1178, 1178, 1179, 1179, 1179, 1179, 1180, 1180, 1180, 1180, 1181, 1181, 1181, 1181, 1182, 1182, 1182, 1182, 1183, 1183, 1183, 1183, 1184, 1184, 1184, 1185, 1185, 1185, 1186, 1186, 1186, 1186, 1187, 1187, 1187, 1187, 1188, 1188, 1188, 1188, 1189, 1189, 1190, 1190, 1190, 1191, 1191, 1191, 1192, 1192, 1192, 1193, 1193, 1193, 1193, 1194, 1194, 1195, 1195, 1195, 1195, 1196, 1196, 1197, 1198, 1198, 1198, 1198, 1199, 1199, 1199, 1200, 1200, 1200, 1200, 1201, 1201, 1201, 1201, 1202, 1203, 1203, 1203, 1203, 1204, 1204, 1204, 1204, 1205, 1205, 1205, 1205, 1206, 1206, 1206, 1206, 1207, 1207, 1208, 1208, 1208, 1208, 1209, 1209, 1209, 1209, 1210, 1210, 1210, 1210, 1211, 1211, 1211, 1211, 1212, 1212, 1212, 1212, 1213, 1213, 1213, 1213, 1214, 1214, 1214, 1214, 1215, 1215, 1215, 1215, 1216, 1216, 1216, 1216, 1217, 1217, 1217, 1218, 1218, 1218, 1219, 1219, 1219, 1219, 1220, 1220, 1220, 1220, 1221, 1221, 1221, 1221, 1222, 1222, 1222, 1222, 1223, 1223, 1223, 1223, 1224, 1224, 1224, 1224, 1225, 1225, 1225, 1225, 1226, 1226, 1227, 1227, 1227, 1227, 1228, 1228, 1228, 1228, 1229, 1229, 1229, 1229, 1230, 1230, 1230, 1230, 1231, 1231, 1232, 1232, 1232, 1232, 1233, 1233, 1233, 1233, 1234, 1234, 1234, 1234, 1235, 1235, 1235, 1235, 1236, 1236, 1236, 1236, 1237, 1237, 1237, 1237, 1238, 1238, 1238, 1239, 1239, 1239, 1239, 1240, 1240, 1240, 1241, 1241, 1241, 1241, 1242, 1242, 1242, 1242, 1243, 1243, 1243, 1243, 1244, 1244, 1244, 1244, 1245, 1245, 1245, 1245, 1246, 1246, 1246, 1247, 1247, 1247, 1247, 1248, 1248, 1248, 1248, 1249, 1249, 1249, 1249, 1250, 1250, 1250, 1250, 1251, 1251, 1251, 1251, 1252, 1252, 1252, 1252, 1253, 1253, 1253, 1253, 1254, 1255, 1255, 1255, 1256, 1256, 1257, 1257, 1257, 1257, 1258, 1258, 1258, 1260, 1260, 1261, 1261, 1262, 1262, 1262, 1263, 1263, 1264, 1265, 1265, 1265, 1266, 1267, 1267, 1268, 1268, 1268, 1269, 1269, 1269, 1269, 1270, 1271, 1271, 1271, 1271, 1272, 1272, 1272, 1272, 1273, 1274, 1274, 1275, 1275, 1275, 1276, 1276, 1276, 1277, 1278, 1278, 1279, 1279, 1279, 1279, 1280, 1280, 1281, 1282, 1282, 1283, 1283, 1283, 1284, 1284, 1284, 1285, 1286, 1286, 1287, 1287, 1287, 1287, 1288, 1288, 1289, 1289, 1289, 1290, 1291, 1291, 1291, 1292, 1292, 1292, 1293, 1293, 1293, 1293, 1294, 1294, 1296, 1297, 1297, 1297, 1298, 1298, 1298, 1298, 1299, 1299, 1299, 1300, 1300, 1300, 1300, 1301, 1301, 1301, 1302, 1302, 1302, 1302, 1303, 1303, 1303, 1303, 1304, 1304, 1304, 1304, 1305, 1305, 1305, 1305, 1306, 1306, 1308, 1309, 1310, 1310, 1310, 1310, 1311, 1311, 1311, 1312, 1312, 1313, 1313, 1313, 1313, 1314, 1314, 1314, 1314, 1315, 1315, 1315, 1315, 1316, 1316, 1316, 1316, 1317, 1317, 1317, 1317, 1318, 1318, 1318, 1318, 1319, 1321, 1322, 1322, 1323, 1323, 1325, 1326, 1326, 1326, 1327, 1327, 1327, 1327, 1328, 1328, 1330, 1330, 1331, 1331, 1332, 1332, 1333, 1333, 1334, 1334, 1335, 1335, 1336, 1336, 1336, 1337, 1337, 1337, 1338, 1338, 1339, 1339, 1339, 1340, 1340, 1341, 1341, 1342, 1342, 1342, 1342, 1343, 1343, 1343, 1343, 1344, 1344, 1345, 1345, 1345, 1346, 1347, 1348, 1348, 1348, 1348, 1349, 1349, 1349, 1349, 1350, 1350, 1350, 1350, 1351, 1351, 1352, 1353, 1354, 1354, 1354, 1355, 1355, 1355, 1355, 1356, 1356, 1356, 1356, 1357, 1357, 1357, 1357, 1358, 1358, 1358, 1358, 1359, 1359, 1359, 1359, 1360, 1360, 1360, 1360, 1361, 1361, 1361, 1361, 1362, 1362, 1362, 1362, 1363, 1363, 1363, 1363, 1364, 1364, 1364, 1364, 1365, 1365, 1365, 1365, 1366, 1366, 1366, 1366, 1367, 1367, 1367, 1368, 1368, 1368, 1369, 1369, 1369, 1369, 1370, 1370, 1370, 1370, 1371, 1371, 1371, 1371, 1372, 1372, 1373, 1373, 1373, 1374, 1374, 1374, 1375, 1375, 1375, 1376, 1376, 1376, 1376, 1377, 1377, 1378, 1378, 1378, 1378, 1379, 1379, 1380, 1381, 1381, 1381, 1381, 1382, 1382, 1382, 1383, 1383, 1383, 1383, 1384, 1384, 1384, 1384, 1385, 1385, 1385, 1386, 1386, 1386, 1386, 1387, 1387, 1387, 1387, 1388, 1388, 1388, 1388, 1389, 1389, 1390, 1390, 1390, 1391, 1392, 1392, 1392, 1393, 1393, 1393, 1393, 1394, 1394, 1394, 1394, 1395, 1395, 1395, 1395, 1396, 1396, 1396, 1396, 1397, 1397, 1397, 1397, 1398, 1398, 1399, 1399, 1399, 1399, 1400, 1400, 1400, 1400, 1401, 1401, 1401, 1401, 1402, 1402, 1402, 1402, 1403, 1403, 1403, 1403, 1404, 1404, 1404, 1404, 1405, 1405, 1405, 1405, 1406, 1406, 1406, 1407, 1407, 1407, 1408, 1408, 1408, 1408, 1409, 1409, 1409, 1409, 1410, 1410, 1410, 1410, 1411, 1411, 1411, 1412, 1412, 1413, 1413, 1413, 1413, 1414, 1414, 1414, 1415, 1415, 1415, 1415, 1416, 1416, 1416, 1416, 1417, 1417, 1417, 1417, 1418, 1418, 1418, 1418, 1419, 1419, 1419, 1419, 1420, 1420, 1420, 1420, 1421, 1421, 1421, 1421, 1422, 1423, 1423, 1423, 1424, 1425, 1425, 1425, 1425, 1426, 1426, 1426, 1426, 1427, 1427, 1427, 1427, 1428, 1428, 1428, 1428, 1429, 1429, 1429, 1429, 1430, 1430, 1430, 1430, 1431, 1431, 1431, 1431, 1432, 1432, 1433, 1433, 1433, 1433, 1434, 1434, 1434, 1434, 1435, 1435, 1435, 1435, 1436, 1436, 1436, 1436, 1437, 1437, 1437, 1437, 1438, 1438, 1438, 1438, 1439, 1439, 1439, 1439, 1440, 1440, 1440, 1440, 1441, 1441, 1441, 1442, 1442, 1442, 1443, 1443, 1443, 1443, 1444, 1444, 1444, 1444, 1445, 1445, 1445, 1445, 1446, 1446, 1447, 1448, 1448, 1448, 1449, 1449, 1449, 1449, 1450, 1450, 1450, 1451, 1451, 1452, 1453, 1453, 1454, 1454, 1454, 1455, 1455, 1455, 1456, 1457, 1458, 1458, 1459, 1459, 1459, 1460, 1460, 1462, 1463, 1463, 1463, 1464, 1464, 1464, 1464, 1465, 1466, 1467, 1467, 1468, 1468, 1468, 1469, 1469, 1470, 1471, 1472, 1472, 1472, 1472, 1473, 1473, 1473, 1474, 1474, 1474, 1474, 1475, 1475, 1475, 1477, 1478, 1478, 1479, 1479, 1479, 1480, 1480, 1480, 1481, 1481, 1482, 1482, 1483, 1483, 1484, 1484, 1484, 1484, 1485, 1485, 1485, 1486, 1486, 1486, 1487, 1487, 1487, 1487, 1488, 1488, 1488, 1488, 1489, 1489, 1489, 1489, 1490, 1490, 1490, 1491, 1491, 1491, 1491, 1492, 1492, 1492, 1492, 1495, 1496, 1496, 1496, 1496, 1497, 1497, 1497, 1497, 1498, 1498, 1498, 1499, 1499, 1499, 1499, 1500, 1500, 1500, 1500, 1501, 1501, 1501, 1501, 1502, 1502, 1502, 1502, 1503, 1503, 1503, 1503, 1504, 1504, 1504, 1505, 1507, 1508, 1508, 1509, 1509, 1510, 1511, 1511, 1512, 1512, 1512, 1513, 1514, 1515, 1515, 1516, 1516, 1517, 1517, 1518, 1518, 1519, 1519, 1520, 1521, 1521, 1521, 1522, 1522, 1522, 1523, 1523, 1523, 1524, 1524, 1525, 1525, 1525, 1526, 1527, 1527, 1527, 1528, 1528, 1528, 1528, 1529, 1529, 1530, 1530, 1530, 1531, 1531, 1531, 1533, 1533, 1533, 1534, 1534, 1534, 1534, 1535, 1535, 1535, 1535, 1536, 1536, 1536, 1537, 1537, 1539, 1540, 1540, 1540, 1540, 1541, 1541, 1541, 1541, 1542, 1542, 1542, 1542, 1543, 1543, 1543, 1543, 1544, 1544, 1544, 1544, 1545, 1545, 1545, 1545, 1546, 1546, 1546, 1546, 1547, 1547, 1547, 1547, 1548, 1548, 1548, 1548, 1549, 1549, 1549, 1549, 1550, 1550, 1550, 1550, 1551, 1551, 1551, 1551, 1552, 1552, 1552, 1552, 1553, 1553, 1553, 1554, 1554, 1554, 1555, 1555, 1555, 1555, 1556, 1556, 1556, 1556, 1557, 1557, 1557, 1557, 1558, 1558, 1559, 1559, 1559, 1560, 1560, 1560, 1561, 1561, 1561, 1562, 1562, 1562, 1562, 1563, 1563, 1564, 1564, 1564, 1564, 1565, 1566, 1566, 1566, 1567, 1567, 1567, 1567, 1568, 1568, 1568, 1569, 1569, 1569, 1569, 1570, 1570, 1570, 1571, 1571, 1571, 1571, 1572, 1572, 1572, 1572, 1573, 1573, 1573, 1573, 1574, 1574, 1574, 1574, 1575, 1576, 1576, 1576, 1577, 1577, 1578, 1578, 1578, 1578, 1579, 1579, 1579, 1579, 1580, 1580, 1580, 1580, 1581, 1581, 1581, 1581, 1582, 1582, 1582, 1582, 1583, 1583, 1583, 1584, 1584, 1584, 1585, 1585, 1585, 1585, 1586, 1586, 1586, 1586, 1587, 1587, 1587, 1587, 1588, 1588, 1588, 1588, 1589, 1589, 1589, 1589, 1590, 1590, 1590, 1590, 1591, 1591, 1591, 1591, 1592, 1592, 1592, 1593, 1593, 1593, 1594, 1594, 1594, 1594, 1595, 1595, 1595, 1595, 1596, 1596, 1596, 1596, 1597, 1597, 1598, 1598, 1598, 1598, 1599, 1599, 1599, 1600, 1600, 1600, 1600, 1601, 1601, 1601, 1602, 1602, 1602, 1602, 1603, 1603, 1603, 1603, 1604, 1604, 1604, 1604, 1605, 1605, 1605, 1605, 1606, 1606, 1606, 1606, 1607, 1607, 1607, 1607, 1608, 1608, 1608, 1608, 1609, 1609, 1610, 1610, 1610, 1611, 1612, 1612, 1612, 1612, 1613, 1613, 1613, 1613, 1614, 1614, 1614, 1614, 1615, 1615, 1615, 1615, 1616, 1616, 1616, 1616, 1617, 1617, 1617, 1617, 1618, 1618, 1619, 1619, 1619, 1619, 1620, 1620, 1620, 1620, 1621, 1621, 1621, 1621, 1622, 1622, 1622, 1622, 1623, 1623, 1623, 1623, 1624, 1624, 1624, 1624, 1625, 1625, 1625, 1625, 1626, 1626, 1626, 1627, 1627, 1627, 1628, 1628, 1628, 1628, 1629, 1629, 1629, 1629, 1630, 1630, 1630, 1630, 1631, 1631, 1632, 1632, 1633, 1633, 1633, 1634, 1634, 1634, 1634, 1635, 1635, 1635, 1635, 1636, 1637, 1637, 1638, 1638, 1639, 1639, 1640, 1640, 1640, 1641, 1642, 1643, 1643, 1643, 1644, 1644, 1645, 1645, 1646, 1647, 1647, 1647, 1648, 1648, 1648, 1648, 1649, 1649, 1649, 1650, 1651, 1652, 1652, 1652, 1653, 1653, 1654, 1654, 1654, 1655, 1656, 1656, 1656, 1656, 1657, 1657, 1657, 1658, 1658, 1658, 1658, 1659, 1659, 1660, 1661, 1662, 1662, 1662, 1663, 1663, 1663, 1664, 1664, 1665, 1665, 1665, 1667, 1667, 1667, 1668, 1668, 1668, 1668, 1669, 1669, 1669, 1670, 1670, 1670, 1671, 1671, 1671, 1671, 1672, 1672, 1672, 1672, 1673, 1673, 1673, 1673, 1674, 1674, 1674, 1675, 1675, 1675, 1675, 1676, 1676, 1676, 1678, 1679, 1680, 1680, 1680, 1680, 1681, 1681, 1681, 1681, 1682, 1682, 1682, 1683, 1683, 1683, 1683, 1684, 1684, 1684, 1684, 1685, 1685, 1685, 1685, 1686, 1686, 1686, 1686, 1687, 1687, 1687, 1687, 1688, 1688, 1688, 1690, 1691, 1692, 1692, 1693, 1693, 1694, 1694, 1695, 1695, 1695, 1695, 1696, 1696, 1697, 1698, 1698, 1699, 1699, 1700, 1700, 1701, 1701, 1702, 1702, 1703, 1703, 1704, 1704, 1704, 1705, 1705, 1705, 1706, 1706, 1706, 1707, 1707, 1708, 1708, 1709, 1709, 1710, 1710, 1710, 1710, 1711, 1711, 1711, 1711, 1712, 1712, 1713, 1713, 1713, 1714, 1715, 1716, 1716, 1716, 1716, 1717, 1717, 1717, 1717, 1718, 1718, 1718, 1718, 1719, 1719, 1720, 1721, 1722, 1722, 1722, 1723, 1725, 1725, 1725, 1726, 1726, 1726, 1726, 1727, 1727, 1727, 1727, 1728, 1728, 1728, 1729, 1729, 1729, 1729, 1730, 1730, 1730, 1730, 1731, 1731, 1735, 1735, 1735, 1735, 1740, 1740, 1741, 1741, 1741, 1741, 1742, 1742, 1742, 1743, 1743, 1743, 1743, 1744, 1744, 1744, 1744, 1745, 1745, 1745, 1746, 1746, 1746, 1746, 1747, 1747, 1747, 1747, 1748, 1748, 1748, 1748, 1749, 1749, 1749, 1749, 1750, 1750, 1750, 1750, 1751, 1751, 1751, 1751, 1752, 1752, 1752, 1752, 1753, 1753, 1753, 1753, 1754, 1754, 1754, 1754, 1755, 1755, 1755, 1755, 1756, 1756, 1756, 1756, 1757, 1757, 1757, 1757, 1758, 1758, 1758, 1758, 1759, 1759, 1759, 1759, 1760, 1760, 1760, 1760, 1761, 1761, 1761, 1761, 1762, 1762, 1762, 1762, 1763, 1763, 1763, 1763, 1764, 1764, 1765, 1765, 1765, 1765, 1766, 1766, 1766, 1766, 1767, 1767, 1767, 1767, 1768, 1768, 1768, 1768, 1769, 1769, 1769, 1769, 1770, 1770, 1770, 1770, 1771, 1771, 1771, 1772, 1772, 1772, 1773, 1773, 1773, 1773, 1774, 1774, 1774, 1774, 1775, 1775, 1775, 1775, 1776, 1776, 1776, 1776, 1777, 1777, 1777, 1777, 1778, 1778, 1778, 1778, 1779, 1779, 1779, 1780, 1780, 1780, 1781, 1781, 1781, 1781, 1782, 1782, 1782, 1782, 1783, 1783, 1784, 1784, 1785, 1785, 1785, 1785, 1786, 1786, 1786, 1787, 1787, 1787, 1788, 1788, 1788, 1789, 1789, 1789, 1790, 1790, 1790, 1790, 1791, 1791, 1791, 1791, 1792, 1792, 1792, 1792, 1793, 1794, 1794, 1794, 1795, 1795, 1795, 1795, 1796, 1796, 1796, 1797, 1797, 1797, 1797, 1798, 1798, 1799, 1799, 1800, 1800, 1800, 1800, 1801, 1801, 1802, 1802, 1802, 1803, 1804, 1804, 1805, 1805, 1805, 1805, 1806, 1807, 1807, 1807, 1808, 1808, 1808, 1809, 1809, 1809, 1810, 1811, 1811, 1811, 1812, 1812, 1812, 1813, 1813, 1813, 1815, 1815, 1815, 1816, 1816, 1816, 1816, 1817, 1817, 1817, 1817, 1818, 1818, 1818, 1818, 1819, 1819, 1820, 1820, 1820, 1821, 1822, 1822, 1822, 1822, 1823, 1823, 1823, 1823, 1824, 1824, 1824, 1824, 1825, 1825, 1825, 1825, 1826, 1826, 1826, 1827, 1827, 1827, 1828, 1828, 1828, 1828, 1829, 1829, 1829, 1829, 1830, 1830, 1830, 1830, 1831, 1831, 1831, 1831, 1832, 1832, 1832, 1832, 1833, 1833, 1833, 1833, 1834, 1834, 1834, 1834, 1835, 1835, 1836, 1836, 1836, 1836, 1837, 1837, 1837, 1837, 1838, 1838, 1838, 1838, 1839, 1839, 1839, 1840, 1840, 1840, 1841, 1841, 1841, 1841, 1842, 1842, 1842, 1843, 1843, 1843, 1843, 1844, 1844, 1844, 1845, 1845, 1845, 1845, 1846, 1846, 1846, 1846, 1847, 1847, 1847, 1847, 1848, 1848, 1848, 1848, 1849, 1849, 1849, 1849, 1850, 1850, 1850, 1850, 1851, 1851, 1851, 1851, 1852, 1853, 1853, 1853, 1854, 1854, 1855, 1855, 1855, 1855, 1856, 1856, 1856, 1856, 1857, 1857, 1857, 1857, 1858, 1858, 1858, 1858, 1859, 1859, 1859, 1859, 1860, 1860, 1860, 1861, 1861, 1861, 1862, 1862, 1862, 1862, 1863, 1863, 1863, 1863, 1864, 1864, 1864, 1864, 1865, 1865, 1865, 1865, 1866, 1866, 1866, 1866, 1867, 1867, 1867, 1867, 1868, 1868, 1868, 1868, 1869, 1869, 1869, 1870, 1870, 1870, 1871, 1871, 1871, 1871, 1872, 1872, 1872, 1872, 1873, 1873, 1873, 1873, 1874, 1874, 1875, 1875, 1876, 1876, 1876, 1877, 1877, 1878, 1878, 1879, 1879, 1879, 1880, 1881, 1881, 1882, 1882, 1882, 1882, 1883, 1883, 1883, 1883, 1884, 1886, 1886, 1887, 1887, 1887, 1888, 1888, 1889, 1890, 1890, 1890, 1891, 1891, 1891, 1892, 1893, 1893, 1894, 1895, 1895, 1895, 1896, 1896, 1896, 1896, 1897, 1897, 1898, 1899, 1899, 1900, 1900, 1900, 1901, 1901, 1902, 1902, 1903, 1903, 1904, 1904, 1904, 1905, 1905, 1906, 1906, 1906, 1906, 1907, 1907, 1907, 1908, 1908, 1909, 1909, 1909, 1909, 1910, 1910, 1910, 1910, 1911, 1911, 1911, 1911, 1912, 1912, 1912, 1913, 1913, 1913, 1913, 1914, 1914, 1914, 1916, 1917, 1917, 1917, 1917, 1918, 1918, 1919, 1919, 1919, 1920, 1920, 1920, 1920, 1921, 1921, 1922, 1922, 1922, 1922, 1923, 1923, 1923, 1923, 1924, 1924, 1924, 1924, 1925, 1925, 1925, 1925, 1926, 1926, 1926, 1926, 1928, 1929, 1929, 1929, 1930, 1930, 1930, 1931, 1931, 1931, 1932, 1932, 1932, 1932, 1933, 1935};

//Conatant array to load the instruction BRAM
localparam integer total_instructions = 2049;
localparam integer sub_instructions = 12;
localparam integer Inst[0:2048][0:11] = '{{0, 0, 0, 0, 0, 0, 1678639104, 0, 41984, -1542569984, 1073741824, 26638},{0, 0, 0, 0, 0, 0, -1542717440, -1073741824, 49157, -1542717348, 0, 0},{0, 0, 1646788608, 14329520, 0, 0, -469762048, 0, 50176, -1475592092, -2140930048, 43022},{0, 0, 1830289408, 18306480, 0, 0, -2079866668, 1088159744, 33805, -603979776, 0, 32768},{0, 0, -1559232512, 15024553, 0, 0, 1685094400, 1073741824, 460806, 1752203264, 0, 25600},{0, 0, -1390411776, 23644552, 0, 0, 344064, 1073741840, 29701, 1946779648, -2147483648, 1049609},{0, 0, 1797783552, 18109872, 0, 0, 0, 1073741831, 458757, -1929347072, -1878523885, 1281029},{0, 0, -1541931008, 13948456, 0, 0, 10587980, 256638992, 661817, 87621632, 16, 0},{0, 0, 1159725056, 13968940, 0, 0, 1342177280, 15, 1453056, 754831280, -810549226, 1004797},{0, 0, -2094530560, 23676341, 0, 0, 0, 116654080, 1028349, -804829452, -2147483633, 1028103},{0, 0, -1541931008, 15021352, 0, 0, 1275068416, 1073741824, 1281286, -49922048, -1068498938, 458040},{0, 0, 1678770176, 19342769, 0, 0, 1688326144, 16, 1049955, 1700986880, 16, 663552},{0, 0, 1259339776, 18262672, 0, 0, 0, -1073741824, 661748, -1265041408, 1330682127, 662779},{0, 0, -1390936064, 18268872, 0, 0, 760905728, -1986789354, 1419526, 755403156, 22, 0},{0, 0, 1243611136, 14002732, 0, 0, -191021056, 9, 0, 10321920, 165150730, 653472},{0, 0, -2062024704, 19350965, 0, 1627389952, 1968887281, 15, 1420639, 0, 1073741824, 1014113},{0, 0, 1244135424, 14330540, 0, 0, -46592176, 15, 1437696, -1862975488, 19, 1438976},{0, 0, -2111307776, 10213941, 0, 0, -2130903040, -1073741819, 360701, 754778112, -1073741808, 1060093},{0, 0, -1574961152, 14374281, 0, 0, 1612300288, 27000842, 1280166, -2002386944, 19, 0},{0, 0, 1159725056, 18142636, 0, 0, 1207959552, -1878482545, 110836, -1331576832, 1, 1050624},{0, 0, 1813512192, 22630833, 0, 0, 2023587840, 22, 1472665, 2013265920, 22, 646297},{0, 0, -1944584192, 14272788, 0, 0, -1543503872, 1437073423, 1438970, -178077696, -1073741803, 1454426},{0, 0, 1679294464, 18129588, 0, 0, -1946157056, 1073741843, 360614, 1554399232, 1197211655, 1281112},{0, 0, -1944584192, 10035636, 0, 0, -1993146368, 19, 1001779, -2013265920, 1073741843, 1002803},{0, 0, -2062548992, 18264393, 0, 0, -1389248512, -1073741815, 634161, -2147483648, 22, 1474866},{0, 0, 1646264320, 10016308, 0, 0, 345590260, 10, 1427456, -1801480760, 9, 661504},{0, 0, 1159725056, 10016300, 0, 0, 1905360896, 421025875, 655671, -2080374784, 5, 655360},{0, 0, 1646788608, 17250005, 0, 0, 1486995456, -1073741805, 1273881, 536870912, 1101004810, 1269047},{0, 0, -1945108480, 20338260, 0, 0, 1499631612, -2147483629, 1420642, 1566248960, 19, 0},{0, 0, -1440219136, 11052556, 0, 0, 288571392, -1073741802, 1258648, 345560624, 22, 1455104},{0, 0, -2094530560, 15423021, 0, 0, 1499091744, 16, 1253376, 939524096, -710410230, 669957},{0, 0, -2094530560, 8865205, 0, 0, 1745520476, -1930422400, 1690331150, -1395719815, -950009856, 60772},{0, 0, -1559232512, 23603881, 0, 889192448, -1474623091, 324009984, -1732196195, 1620902320, -2147483648, 24588},{0, 67108960, 1956270976, 816528691, 1715775625, 915422506, 1813305629, -2131225408, 260089356, -435388304, -1189005632, 58886},{342016, 67, 1952055296, 1903778293, 2082787401, -1727519960, -1039507328, 545785856, 1589665292, -2012348151, -1779656448, 57360},{0, 70778960, 24576, 12298944, 1766651136, 647242654, 1822786156, -2029250176, 1891681798, 1711972460, -1046698560, 60016},{276480, 80, 24576, -1653228224, 1797303625, 160185510, -704094088, -2141714048, 729865735, 1493717861, 1387790336, 33590},{327680, 117440579, -1744830464, 1701555882, 1277480777, 215038888, 168137621, -1341288057, 960521840, 1778749453, -1073741824, 1102225},{327680, 67108976, 24576, -1326106336, 1498191721, -1575928424, 1463373652, 1330471552, -184518855, -1695184348, -701759488, 1050368},{458752, 70254592, 20480, 278495232, 1228723897, -817025700, 50206260, 1345585159, 1666596047, 188280665, -1880816752, 23285},{274432, 117440592, 0, 11124288, 2086456832, -1923734702, 1319219125, -1881839665, 1741918727, 107974613, -2147483632, 457101},{0, 69730416, 24576, 12148256, 2067855360, 55913118, -66775643, 275579718, 1519791621, -1291979883, 275513359, 1005168},{469762048, 67, 20480, -258224672, 1547227825, 533346, 1889617756, 800260432, -205064451, 1889634144, -804457520, 31494},{0, 117440579, 20480, 628735680, 1522063441, -1575732638, -1265004716, -281250353, -1718589640, -17068112, -950271994, 21235},{-2147024896, 66, -1476370432, 1895152333, 1546712217, -1924579820, 1721339121, 1771658000, -1919536384, 888343793, 1251537686, 664411},{0, 70254592, 21376, -248166112, 1255717049, -1546357922, -123858888, 272147401, 738843948, -1829017083, -369319863, 1004193},{-2147076096, 66, 1476395008, 16505293, 2083035136, 1729311320, -1419577835, -1350738027, 628486, 2103433360, -1735301297, 1448287},{0, 70254592, 2013287296, 1903811153, 1732286633, -1542178154, -43706980, 362587157, 1607701861, -627036139, -1340541559, 645791},{339968, 0, 17280, 1891350848, 1143255913, 51133612, -212144159, -1892590955, 1060952, -715472896, -1517751537, 1447671},{327680, 67108864, -2013240448, -377890219, 1546426489, -1496436064, -1843702884, -1026544429, 436550681, 1453770044, 1639266767, 1049439},{342016, 100663360, 0, -489043616, 1279317841, -166973908, -765976140, 1352480015, 1498406427, 788580741, 1233475920, 1007925},{-2147211264, 99, 1879048192, 1865006640, 2067060841, 1745495382, -1633279767, -1189567551, -1849007304, -1466329467, -1058495488, 27658},{-2147090432, 67108947, -1744830464, 16103753, 1808324608, 1699556880, 1265569821, 543165519, 1666189851, 504139693, 374865930, 1027330},{-2147090432, 50331715, 20480, -591806904, -1590388551, 1481203820, 2047255948, -1435982314, 1481216871, -281459316, -2054684672, 646822},{-2147084288, 112, 17024, 816555730, 1732032681, 891024, -1509117128, -522122801, 181794314, 1644712761, 546126272, 1421155},{-2147020800, 83886144, 24576, -1384677376, 2083051633, 1892261018, -1911234456, -1448004973, -1693817329, 1577531216, 321650695, 362357},{340032, 35127296, 268452736, -556750830, 1530435737, -1618266596, 859349122, -2147483629, 4229785, -502222715, -526645824, 1259252},{342080, 101711872, 268451840, -1676997545, 1548520009, -1844495194, 513466483, 412352531, -1991011015, -2106525403, -805003178, 1254144},{-1945763712, 83886144, 28672, 10562592, 1818015744, 1406041634, -1777885030, -1333315767, 1427973, -80001732, -1890278839, 662261},{-2147143680, 67, 12288, 1562869760, 288159929, 1527337057, 456597595, 909468441, -821721440, -452897220, 217317391, 1102692},{65536, 101711872, 17052, -243859456, 1816967273, -1710665706, 251483668, 1404147216, -1777927837, 581071793, 1935579658, 107319},{331776, 70369280, 0, -1331187712, 1278781881, 1167235162, 727968313, 265289750, 1880381706, 56308574, 1245539152, 1041925},{-2006581248, 117440592, 268451840, -1523073003, 2083305329, 332473900, 929350012, -271123533, 109678087, 376420008, 25258646, 1455973},{264192, 1191182384, 21248, 787489824, 1965865089, 739350060, 570766337, -1986782381, 1076889, 984355520, -419219030, 1420037},{-2147479552, 85459043, 16512, 1543503872, 1423493721, 1524071978, 1862743473, 969149008, -1673430321, 1325513141, 548405270, 484097},{201599360, 113, 0, 1903624192, 1817745513, -1643016090, 1385750962, -1440309165, -1614163211, -1164031528, 1331754191, 1440095},{0, 33554432, 17028, 1677721600, 1882765433, 92970541, 2091237832, -1067911153, -132778843, -1688234472, 909780810, 1273746},{262144, 84443136, 384, 15748128, -425641984, 139091502, -1825865464, -2147483639, 5248016, -291477021, 1925007381, 655006},{-2147221504, 1, 58872580, 825744980, 1524160601, 248348834, 1871845672, -271296446, 240090975, -1986871056, -166003131, 679449},{137216, 69746688, 0, 805306368, -262895015, -1919828576, 1533013845, 328038287, 968995867, -1154059365, 18, 1629184},{131072, 0, 16384, 436798816, 836016305, -1814594663, 865472385, 272733136, -133367601, 1627642208, 217908303, 1646325},{196608, 83886112, 16384, 814448640, 551073945, -1752135649, 1869256928, -656670710, 1795845642, 1376704129, 1491113935, 1453928},{327680, 1048576, 1879064576, 393861621, 355768465, 1812744289, -166948803, -1874762484, 831499611, 319434813, 1448423824, 1063787},{0, 80, 16520, 817607729, 1472760497, 1703506154, 1626605945, 1244226951, -1747550554, -1364818076, -375458752, 1628686},{262144, 84459521, 67239936, 821406325, 1260697489, -200200676, 926109852, -1288145392, -180303005, -1426393354, 21, 0},{137216, 69828624, 0, 393854656, 1464391849, -716339160, -1973884496, 1291423173, -212624653, 1047931418, 15, 0},{-2147483648, 66, 256, 805306368, -237193063, 798140524, -995862243, -221993838, 483059, 1167201020, -369279094, 1286963},{329728, 70303744, 8192, 1902116864, 1548523705, 1733244004, -214781939, 1405434060, 965325671, -621594797, -1877893800, 1257273},{272384, 16777312, 1342177280, 820754114, 1252841625, -174967528, 1057206406, -1969159862, -1441611019, -1620699448, 9, 1049600},{69632, 85458944, 63062016, 23077930, 1269610496, 1536335394, -1767868883, -700884205, -745533597, -1819119820, -1925709800, 1472355},{272768, 48, 4352, 621829120, 1815656569, 1410549274, 1129969234, 29201994, -1772898663, 1520043333, -1239934129, 666423},{-2147477504, 67108944, 0, 821371922, 1278785721, 961654950, 928739377, -1286260330, 1502556929, -1364997751, -1968372907, 624985},{201326592, 83886147, 0, 1899464000, 1549586065, -1836218218, 974657825, -206396266, -1878863277, -1553659323, 1, 675216},{4288, 69730304, 134242432, 1899736781, 1462013777, 173159952, -1553238949, 1337785104, 38806794, -1768396387, -375587883, 1267363},{0, 1157677056, 268452612, 1895085109, 1548519609, 1770923564, -1267661055, -690920683, 1506218338, 504673962, -162392007, 672262},{0, 1627390048, 17032, 10500096, 1480898304, 223059102, -1709948608, 14155785, 226517516, -1173323572, 872852705, 1465090},{-2147221504, 33, 4096, 826310656, 474142073, -1605198289, -2039443076, 1900871877, -1604733028, -1290268656, 1247876288, 1422961},{131072, 67633248, 20480, 704643072, 473209009, 248495261, -100019524, -1050855147, 734061065, -2036440755, 1625635776, 36598},{395264, 68157520, 134230016, 1702345322, 1549323613, -1987465684, 245753225, -1445199865, -1996026017, 1847408793, -1981768320, 162713},{0, 1124073472, 17028, 1693538368, -1404791439, -1584685522, 173279784, 218156801, 117468166, -2112123048, -266654732, 40453},{-2013265920, 1572928, 0, 23101440, -1255892992, 332299748, -120631980, -1188638836, 1410897496, -208474788, -2059403264, 81926},{262208, 0, 12288, 818940352, 2084712361, 168992301, 1041986463, -1987774395, 1087894, 420024196, 426285127, 1542769},{0, 83886080, 16652, 485818368, 1355585713, 1526313, 1661173924, 20710863, 332413963, -428767472, 809896719, 849668},{-2147090432, 524354, 8576, 590825824, 1750915153, 118041370, -703807296, -1246756849, 114909807, -2023022388, 1618041558, 1631118},{4288, 67108864, 20480, 0, 1757585664, -49308521, -1083428798, 1409577109, 1089836, 40976384, -738692793, 22323},{131072, 16777216, 12288, 0, -71641856, 1203732, 773144788, 22547914, -83203570, 1712308568, -2124874809, 1000975},{262144, 33554480, 0, 613416960, 1891932241, -1542743199, -1020024184, 1073741842, -79206748, 1185042360, 1243675535, 693410},{0, 17874944, 0, 1509949440, 961989196, 1665891869, -1117809095, -2094964861, 349124344, -7459494, -2141701236, 1472760},{6144, 68157520, 0, -1040187392, -1495758707, -1584694382, -962289328, 1450704914, 1829373452, -12601639, 1249994889, 1453077},{340032, 118489152, 134217728, -1452550552, 1221154906, 164572690, 1526199927, 1364721664, 210731763, 463302801, 1330443606, 1297243},{-2147481600, 33, 0, 469762048, 2086283642, 1879807509, 392569268, 654640720, 118934186, -1314781435, 25, 1683874},{0, 80, 16396, -1340831200, 1279088786, -1734910436, 1838436236, 25, -1559239005, 1838436236, 902010521, 1039204},{6144, 33554432, 16384, 437977088, 2032176201, -1748001251, -1575214772, -1784820151, 63658, 1190419684, 256203269, 1629848},{272768, 558592, 0, 1830280224, 1781831025, 831206936, 1056455011, 25, -1427051277, 1519957402, -897539629, 1252709},{-2147418112, 83886177, 1342193672, 825699917, 1818003849, 1653616172, 661231149, -157195175, 1681960850, -278066459, -1437637888, 622244},{67506176, 67108976, 20480, 1879048192, -1134786487, 277909012, -888512296, -265945088, -36720901, 456774540, -1052439981, 1463816},{262272, 83886128, 4096, 1899462656, -1187579791, -187320790, 1533880082, -798409642, 952476422, 2131152737, 1101004809, 1482267},{-2147483648, 0, 0, 1197473792, -329440686, 1468759578, -1196911684, -209090349, -2000627188, -1254767235, -1068214317, 40980},{-2147221504, 33554433, 4096, -1577058304, -63244180, 998856230, -1298280311, -268093303, 464660, -2096611328, -792920047, 1147549},{131072, 69730400, -1174138880, 1832368875, 743757923, -892776215, -1620568456, -1934884864, -1563820382, -7195714, 7119250, 61959},{262144, 118489088, 21248, 0, 724137984, -740997029, 260683472, 16, -736740352, -1684427524, 544039699, 1284865},{-2147155968, 65, 4096, 24707072, 1814381056, 1783716843, 1523593085, 1888323855, -741385644, 275781992, 222035975, 667529},{0, 68681824, 20484, -1327462368, -1134784591, 22048, -1923377752, -741786541, 970340874, 987095217, 754910221, 1456660},{-2147483648, 66, 8192, 116739360, 1625077873, 813093, -936568660, -1597142336, 760833889, -1450157668, 1493445974, 1093467},{131072, 100663360, 20480, 615579648, 280926365, -1730824675, 1047580832, -114294768, -1827431917, 1041170669, -1985999094, 1062653},{395264, 69730304, -1475215360, 821746283, 1546161521, 13803672, -2113458155, -851967999, 1937826195, 56964529, -1723804775, 1508609},{0, 83918896, 16384, -249069568, 1549345109, 1477145409, -1324855284, -1977284535, 1490290427, -1636732214, -1970756471, 630434},{262144, 1572880, 8192, -1322931680, 203544699, -1508459965, -1230419572, 1250208341, -1690215672, -1106253284, 174627663, 88744},{196608, 524288, 180748288, 17844265, 1789559296, 1087356455, 1175230073, 1286417674, 1476776, -1163761124, 212938063, 1476776},{268288, 83886096, 24832, -1493860352, 1545982637, -49627614, 104591560, 266665418, 114264841, 303423816, 1902384144, 680498},{327680, 67126784, 8192, 12167744, 1750898688, 952282641, -1099939408, 1073741842, 1839321095, -1083659645, 1081618450, 87580},{262144, 0, 0, -973078528, 551215700, -1857324125, -1954589291, 1192521925, -1726501505, -1401861728, 1494745111, 1090393},{-2147483648, 68206592, 20480, -1320124416, -1473324870, 626194, -1196697356, 1789433866, -1747946896, -1147454942, -1957851263, 1007256},{2182, 67108864, 0, 715905312, 959484041, -118587877, 1805056326, 1120927769, 1260590, 1127338233, 1396781893, 1489249},{-2147477504, 66, 4352, 1891322944, -95111087, -1576456668, -89475376, 1983483136, 1017496, 495779840, 916284298, 86680},{0, 16, 8576, -1060044800, -1256114061, 1152544, 358400000, 365494672, 1560970043, 425512977, 806444240, 1253222},{0, 50331648, 0, -986284032, -1339407950, -1449695724, 1813730876, 16, -183700480, -147222688, -1980182646, 1458531},{196608, 17, 16384, 821723136, 651250825, -971737897, 1184909157, 1012924417, 1976802833, -1489251400, -1970456752, 1261369},{-2147418112, 33, -1476395008, -256356256, -1811564429, -1856547284, -949087359, -259704813, 1008390, -513550056, -694328503, 1053026},{0, 0, 0, -948371456, -1867865486, 756448794, 1889702813, 329067776, -29270521, -2059824988, -1818162474, 662841},{272512, 0, 24576, -252978580, -1675061078, 1674723418, 996126911, 372830998, 80902, -1667232056, 824503434, 1473182},{0, 33554432, 274202624, 24757332, -716622166, -166823196, -1919515844, 257492496, 101690614, 1915978145, 0, 1072128},{327680, 33554480, 16384, -253394944, 274612564, 797732385, 906695621, -1818412657, 1496923, 1130089012, -1976225843, 1424218},{201326592, 65, 0, -1387167744, 735183211, -1890630429, 1228378953, 963336733, -1887323285, 453758985, 1400714439, 53528},{-2147155968, 64, 0, 482071584, 828007249, 1603357541, -1963616771, 552689609, 668171, 621514676, 320932755, 1425162},{-2147483648, 101711937, -1442819968, 821800650, 1545918625, 882214, -815032572, -155618176, 1633478553, 1200649801, 910779791, 1418091},{65536, 0, 12288, 1159725056, -1404111283, -1991543976, 385188253, 123739079, 656630, -227157868, -815499712, 632488},{65536, 64, 0, -973078528, 1255793306, 1745494948, 1520961940, -1982794367, 1750484646, 1016942752, -1982526966, 1055401},{264192, 0, 0, 91684864, -708400564, 1473492516, -620207968, 92109952, -960131574, -936535752, -1724332329, 360493},{0, 0, 4096, -2030337504, 651526733, 483105685, -1389210852, 1493434389, -1874743141, -1254991579, 1495309142, 1085330},{-2147483648, 83886144, 1207985032, -1493845683, 1808312417, 877739428, -870642507, -1397212799, 1609576, 2115333300, 873673861, 359946},{65536, 0, 8576, 824690016, 204920165, 856249263, -1701245711, -863764464, -934477517, 1248954784, 1829031745, 1103639},{266240, 0, 0, 1186693120, 1263048861, -824924068, -1372571488, -856948724, -1685486200, -963077992, 433363841, 699786},{71499776, 67108944, 0, -249056224, 1547881090, 361872925, -166772520, 655850231, -1421017446, -10387204, 12, 88226},{0, 68206672, 1744830464, 1895161408, 10892881, -967954927, -442836671, -642935806, -1571253715, 1051519850, -2147483635, 187846},{0, 1048624, 16512, 1879048192, 1809239571, 923749905, -1940352139, -980601019, 999358300, -278152907, 806982466, 1065780},{327680, 70795296, 2013290880, 1788598880, 1280366737, 537680, -1361850520, 222623384, -1613323530, -681871714, 1868354626, 186221},{196608, 16777280, 1342177280, 472204320, 2068493401, 1557118503, -1287941239, -1671352493, 794374969, -827845699, -1781414315, 701601},{0, 33554496, 20484, 627671040, -1579902887, 1782611490, 1029933497, 22, 1636645376, -895756623, -163406829, 1655465},{-2080374784, 33554498, -1207934080, 1899474506, 1815754818, 1421530, 1543503872, 1941908947, 902806178, -1765059879, -1486148086, 666276},{4096, 68681728, 0, 805306368, 1356369241, 1012366249, -1955973651, 1558446096, 1590692303, -1217482443, 331954569, 1458527},{131072, 50331648, 17024, 370212864, 1547212953, -1454080486, -1626992496, -809985837, 47223035, 788418493, 816777546, 1234635},{0, 16777216, 0, 103022592, -1252398732, 1821480494, -1188049744, 1459669781, 695971, 1114406912, -1716178943, 1420633},{264384, 0, 0, 1162870784, -172338813, 202874412, 116794175, 254909447, 1435525899, -1046325068, 1488213401, 1053090},{327680, 18350112, -1404682240, 1903614571, 1546164369, -967557102, -1760702644, -809983403, -963392771, -1566348756, 279225043, 1645408},{0, 33554512, 16524, 452311360, 732992329, -1568651741, 342951684, -162985209, -217480437, -2020783588, 2102365521, 1637210},{131072, 67108864, 4096, -1325685696, 925508356, 39171607, -17430687, 1073741845, 466999554, 520856000, 27090387, 1256054},{201392128, 65, 0, 455081984, -329853863, 1277486, -1160806400, 928423254, -652684431, 1243349436, 27056342, 689318},{0, 67108864, 384, 24677024, -1866429696, -967879764, 1774656912, 28, -960495616, -746814083, 1621411477, 115369},{327680, 524336, 17152, 19955712, 1277988608, -1685567318, 1865554213, 1495611472, 698162, -1566739580, -1246127280, 850459},{262208, 48, 134217728, -1329879038, 1280874603, 764683242, 1644832127, -1733033956, -107492661, 1074238168, 414513537, 834763},{327680, 70254640, 4096, 790648832, 1502435417, 143763612, -2100293939, -855847213, -808012052, 446576934, -1875587303, 119560},{-2147209148, 50331731, 0, 1358285120, 1815648138, -877908454, -771281738, 1641253138, 461402984, -1633576800, 278984131, 701468},{0, 67633152, 0, -2034663424, -247163220, -1995876886, 1060131741, 419430419, 973124912, -895852363, 1485934606, 86320},{262144, 48, 0, -1006632960, -64904844, 936009234, 1779241805, 323827673, -1952852467, 1411258501, 411405185, 1613342},{-2147153920, 33554433, -1342160896, 824565071, 1547995561, 126757904, -1307205384, 959710976, 126531436, -32550024, 1400396032, 1244687},{71680, 1140850688, 1207980828, -1359627955, 2085140121, 118570328, -543494304, -905603582, -1765613911, -99319487, -523096392, 1265463},{69632, 50331712, 461504512, 10529874, 1188599808, -1706058286, 1985541009, -1431002541, 717288251, 933332568, -2041042215, 1293721},{-2147483648, 33, 0, 1769472, 1992704000, 1473224221, 1896272620, 1720518416, 1477264084, -2002892320, 166014726, 1458281},{264192, 0, 8192, 821410112, 832870249, 759738405, -1767343815, -757830504, 1821143448, 1905839544, -843579380, 1295251},{327680, 67143168, 1073741824, 318484161, 1513134225, 1560965991, 1788580593, -755933942, -1674985063, -2023020098, -910074554, 1676696},{0, 69828608, 4364, 490200640, 1211412817, -1986647464, -1120578735, -1735131121, 909333897, 1871946459, -220003508, 834349},{-2147477504, 66, -1879043840, 817487478, 1546170505, 46735914, -149674175, 1830052124, -782694757, -1258121832, 901538133, 1297247},{201326592, 1, 16512, 21037056, 1787131904, -833514015, -2001253099, -258280499, 695035, 80829668, 1890889803, 1264393},{137216, 83886144, 1879048192, 1891224033, -1070286663, -174707180, -1217318692, 1451845721, 1594656510, 453662345, 7, 1003871},{327680, 68681825, 0, 427252128, 1549064281, 97163368, -274559252, 655665996, 97094556, -1146982672, -581590327, 1098402},{0, 16777264, 0, -252411904, 291051525, -2020696933, -980248295, -949685296, 1096219, 779507836, 282132746, 1106458},{339968, 50331648, -1879031808, 1467464386, 1814599849, 277426278, 1117941939, 1351943833, 155877538, -688452991, -814673704, 1862351},{0, 67108947, 134222080, -252988366, -1876330332, -829049310, -708408051, -1244017003, 1429249, 459100920, -218574576, 485213},{262144, 33554432, 0, 370442240, 405310905, -1500537699, 1798851180, -912239665, -1714780506, -1818535648, 1162346509, 1255578},{196608, 1073741888, 21252, 494513856, 1817491537, 1519203620, -895936783, 29890455, -1718421693, 1865793992, 1014487420, 1861469},{0, 33554448, 0, -2038410208, -188287381, -859136476, 654855404, -803681069, 1796441948, -956199679, 1351404822, 971114},{131072, 0, 16524, 1879048192, 1547334283, 1490463, -627435840, -1985959534, 1526809240, -1398171979, -323053110, 1286663},{131072, 50331712, 268435456, -2101748120, 399876213, 1834324627, -818932988, -2102657010, 1834369637, 120623868, 106441421, 47213},{262336, 16, 0, 1140850688, -1177979548, 1435401626, 1661663394, 379365968, 115562, 1353288092, 327177686, 54581},{272384, 16777328, 24960, 791004488, -425420679, 743780524, -892654167, 1626605510, 1208628747, 1395413693, -1602435327, 1246000},{4288, 69730320, 402653184, 8397898, -925070592, 1804432612, -751504513, -2147483648, 1015109490, 1535866661, 427921861, 1296698},{0, 67633152, 20736, 824223763, -341010255, -716212710, 2064274268, 0, 965537792, 1779397565, -211733044, 1442319},{0, 17825856, 0, 570425344, -1747150735, -196452848, 1024150228, -370865325, 1905675158, 1252682128, 322762625, 1078580},{264320, 48, 20480, 805306368, -1254498135, 286754348, 648772006, 1293418512, -778422387, 227793108, -1938765951, 1009242},{65536, 64, 8576, -1837053952, -330467934, -1999143380, 1928060005, 1505074256, -2000037992, -409871255, 964750345, 429673},{0, 50331680, 17048, 824690125, 1814593881, -1572065838, -1651798076, -809195441, 1675001, -1154119040, 1703121901, 813578},{-2012938240, 50331712, -1476395008, 1903672011, 1548523673, -980784028, 648205000, -373103911, -975624549, -1496314432, -903271207, 1676962},{2048, 68157520, 0, 751861760, 1247066257, -212943646, -1690996560, 1102678104, 488158877, -1693865336, 28936271, 693277},{0, 18350081, 16384, 821800640, 1278777497, 611674, -2010316800, -279433898, -1987623166, -1090293599, 1356959829, 848630},{0, 50331664, 8192, -1053458432, -1480972107, 1628018194, -1124023968, -1050648304, -2003988725, 111329769, -1735812405, 752158},{327680, 102236224, 0, 825937920, 557627481, 936021, -1839653796, -1517266280, -971439256, -1559337559, -1817888941, 114715},{0, 69829632, 1744834944, 1903811136, 1730719577, 1532079378, 1835013565, 50605328, -714116768, -1148689949, -167683112, 703394},{0, 119013473, 17024, -251985920, 1522053970, -1698150300, 1546324652, 855157446, 727267085, 2064475744, 959342163, 1276505},{-2147483648, 68157440, 12288, 822149120, 2068141317, -862806505, 1030968725, 625572997, 1087144, 1727478988, 88688783, 1117863},{2048, 69779488, 0, 1898020864, 1465159513, 403946920, -681727592, 21, 1834774125, -1369066758, 364731266, 446812},{397504, 67108864, 20608, 820749376, 1549195417, 101360790, 1118239163, 22, -799455232, -2108379000, 2035127301, 1241754},{333824, 65, 0, 807075840, 2082509177, 894065221, -683429019, -1346303086, 910608924, -1062516191, -1822949361, 1505078},{339968, 16777216, 16396, 15826944, 1895825408, 1800428189, -751884771, 1073741845, 1531780459, -1302213343, -318320170, 1431304},{262272, 16, 0, -2035580928, 1229756523, -1449756072, -1083430494, 90033871, 663395172, -1667264779, 1383596054, 859375},{397504, 16777296, 16384, 1879048192, 1479841393, 735149526, -1704122665, 21, -1425205760, 187470976, 1789959635, 399152},{272384, 0, 268443648, 821377330, -803161959, 46958702, -422484159, -1940838500, -25002754, 687702652, 1383596048, 351941},{69632, 68681728, 0, 13664256, -1216348160, 1984871956, -960026776, -2023934446, 907313979, -220534935, -2147483627, 485687},{201601024, 84410369, 2082209792, -1321916847, 1818024041, -1386858984, 1584492412, 1999280384, -1713798292, -214125760, -2147483634, 892111},{0, 69730400, 140, 15780896, 1464148480, 1679267216, 281482913, -588984051, 485326, 2121692828, 817090328, 875318},{266240, 0, 4480, 1893826560, 1007024194, 977450543, -16026711, 12, 461492224, 1335646496, 567382607, 711476},{262208, 50331680, 20480, 22085632, 2068624384, -1710124323, -367974998, 1447034908, 1594651501, 2070615717, 161836364, 856826},{331776, 0, 16524, -1342177280, -128141717, 751531540, -2019791664, 225455315, 1672909, 752451584, -1177888374, 1256347},{71680, 1, 0, 11248672, -159383552, 1481348188, -1627622548, -210982705, -1551202421, 5802636, -980680688, 1097014},{333824, 33554448, 17152, 1534689664, 1279834201, 1708207522, -823936872, 1119382732, 1825375846, -971695868, 644098957, 840429},{0, 16777216, 256, 100663296, 1967732291, -930186021, -1989405260, 32074584, 87357, -750941044, 1934182657, 120489},{-2147483648, 524354, 1879072768, 624396995, 1546170713, 865838, -1853256624, -1589590765, 1497542245, -1358028348, -743863856, 47631},{0, 17874944, 268452504, 15452212, -1498589184, -195840670, -1096235244, 274464784, 1615488257, -343361105, 864200961, 55093},{134283264, 67, 134238208, 124366511, 1815656533, 847848996, -1835335407, -441839419, 62983, -1023572200, -1825754495, 32267},{69824, 0, 0, 384892928, 1816582316, 122861103, -1084215145, 1240490325, 1632662900, -392229720, -1774925175, 200350},{0, 17874944, 0, 1879048192, -1253231099, -1915914706, -1351837415, -2147483638, 1540984156, 1647011431, 417435078, 1494424},{0, 16777296, 16768, 1698150752, 1447379561, 1783637458, -1056074308, -1363079794, 648788, -1554266460, -59930092, 1079164},{-2006908928, 100663362, 0, -1341685760, 1817585793, 739728019, -755231667, 1725066593, 1745689485, 1060542125, -971480743, 1299818},{264192, 83886080, 24576, -1418241632, 1546426521, -976079596, -1895255348, 331127960, -1668101100, 1779733408, -528663524, 967572},{137216, 67108880, 0, -246369280, -148858699, 679442, -1163155356, -691183792, -2037398881, 1537513164, 377006547, 1272682},{-2147479552, 67108881, 20480, 825720832, -1497319751, 1746039522, -1235096364, 915156822, 797777618, 1600702944, -858232756, 1232429},{131072, 50331712, 0, 821755904, -1607589527, -1706124142, 506534008, 1175990541, 1607284, -233404900, -1736664420, 92257},{327680, 16777280, 0, 515615424, -333145959, -980603774, -1948970860, 867989142, 186186, -1277820928, -1871395382, 1286614},{-1945884672, 96, 256, 1790683857, 1228445849, 231222098, 303444197, -1344586426, 667394, 1362973540, 718838223, 476931},{0, 67633152, 0, 817613856, -2125165239, 995513892, 1808719081, 7, 1112845312, 1651946537, -1821558884, 857403},{0, 1097792, 0, 0, -374775552, -287873638, 1909250392, 8206922, 474968743, -1028788830, -823132144, 1278357},{69632, 64, 0, 478216192, -1529429895, -976200146, -1563348803, 1249944278, 26409640, -1727115039, 476053514, 1008908},{0, 68681728, 20480, 816555712, 550306473, 1506880799, -1053682271, -710934509, 1020512572, -811797731, -1382494948, 684946},{0, 16777280, 0, 816545792, -2033553055, 1473116, 872415232, 1703477383, -204890259, -1297887044, 1354003350, 1274176},{4096, 68681728, 0, -267386880, 1490145362, 68337055, -757651607, 1343266956, -1602136970, 114927384, -1874525171, 54390},{131072, 0, -1879031808, 817504321, -600153271, 1544191488, 1866273405, 1384209427, 691802, 335544320, -1823450410, 1268587},{201326592, 17, 0, 20414464, -1255786878, -15567314, 757860116, 1656422164, 721838694, -59664092, -651678976, 1315071},{0, 69730400, 8192, 628719616, -1597715535, -863412182, 1758271653, -1031486134, 675634949, 2062509848, 1487523026, 1352397},{65536, 67108896, 1880633344, 1895161450, 1814075557, 618003, 1241513984, 1334376513, -125712581, -885861540, 13977170, 1289745},{469766144, 67, -1476374388, 1891347145, -331550055, -1912363486, 1593914289, -1568760176, -1995277570, -443705183, -1433204840, 808692},{0, 68681808, 4096, -1328513024, -1589331877, -1768973166, -544237203, -864446769, -963419300, 1655421152, -1728213101, 1257159},{4096, 67633200, 0, 11553824, -698836992, 1695448622, 2004186717, 16, 1409938090, 1117693252, 1448912019, 967764},{268288, 16777216, 256, -455081984, -1257621429, -1722565206, 1939417828, 476120268, 1475910, -2084155316, -350407335, 1631084},{2240, 0, 8192, 8388608, 2066083328, 810638869, -1010372390, 1138253198, 901964848, -802257960, -1073741806, 1615453},{0, 16777248, 17024, -952682944, 2083190922, 1568769581, 459245332, 98129222, -1852581216, -1364600231, 796218710, 632570},{272512, 18350080, 0, 815378496, 1270387321, 1758471010, -828181809, 1200096130, 1850336366, 1254504856, -947125375, 1295256},{-2147483648, 0, 0, -952771008, 285390963, -930433509, -1805788848, 747644044, 383176554, 1086953900, 1284243458, 385429},{-2144993280, 50331714, 8192, 590719575, 1815656569, 99858, 108085248, -158422215, -557396087, -86500248, 1307377154, 189397},{-2012866560, 67108944, -1413480448, -1330927928, 1506839921, 873604632, -1976486067, -1507891240, 1904339553, -1911114944, -750454964, 1106165},{264192, 100663344, 20480, 503316480, 1277542993, -1563709926, 1396435588, 49582988, -820153688, -1756703903, -1563126843, 1613577},{0, 68157456, 0, -268435456, -450813772, -2041872850, -1463007352, -1933281140, -493627572, 112047304, -836204906, 685258},{0, 50331648, 4352, 12172352, 2067120128, -1810737629, -247735995, -1723596778, -1831619182, 727372641, 922587540, 1293263},{-2147479552, 85459008, 0, 1790696040, 1219014545, 1901341276, 1933227444, 796393482, 1514542621, -1412615263, -1784320180, 1296690},{0, 16777248, 16396, 1409286144, -1212033629, 1228194, -2133655552, 1453642511, 1615497021, -420194639, 715847824, 1426188},{272384, 50331664, 0, -1331676160, -519751587, 1901248016, -1487145566, 482344966, -1663840510, -1502179260, -1877095347, 642309},{264192, 83935232, 0, 1901690880, -150887799, -968120796, -1029103168, 28886671, 1804998791, 1795912711, -2005656557, 1299765},{0, 64, 134222208, 515443118, 2082928705, 1750187541, 449676936, -964352048, 641640, -1993883648, -321071290, 1066517},{0, 67108912, 8192, 356220928, 2171273, 491492767, 1546149056, 30698064, 1213388, 1785824932, 266405256, 372391},{-2147483648, 17825793, 17024, 1899421248, 1262786649, 1387160, 1557664484, -520802740, 1993343811, -12492528, -1486043633, 427725},{0, 97, -1924906356, -2093523370, -600983391, -1967108588, -1862528839, 1889110808, -1962457560, -1819668287, -329578230, 633735},{134217728, 80, 16768, 828997632, 1473285033, -888237996, 1896533172, -1279079604, -163091720, -54030176, -110100456, 810822},{0, 16777216, 8192, 805306368, 1462678125, 1636809965, 1502990073, 1448973782, 60334676, -412133964, 1077502424, 1292143},{4096, 0, 16512, 10498080, -88702208, -720126564, 1869444745, -1979599911, -1277398866, 1952827285, -430147236, 857999},{0, 33554432, 268452480, 817610065, 1087157681, 684290917, -1574024904, 154675402, 876759, 1177374200, -310326011, 979861},{196608, 0, 1342193920, 825735533, 1179009465, 46624, 1851116756, -895978540, -845762984, -1871461024, -1448779771, 1860275},{65536, 67108896, 12288, -243672512, 1279617650, 1402912, 117295420, -1881639869, -1299981646, -694105364, -890465268, 221856},{131072, 48, 17048, 653998752, -1601603479, -1747897564, -814622868, 1466783126, 1436183388, 2002536829, 630157839, 473911},{-2147483648, 16777281, 8192, 582680576, 1185451641, 1645387090, -1290846147, 2032665546, -7730578, -1752065664, -1862704551, 1682175},{262144, 1048592, 12288, 758611968, 1221888913, -686328294, -1026122548, 1298166165, -146650508, -1765166268, 119275532, 1687501},{-2147155968, 67143280, 24576, 1421597280, 1814343593, -1814925796, -214772767, 870421647, -555680040, -1291960990, 330905346, 1649459},{131072, 587202560, 17048, -1331054560, 1792575929, 1817151524, -419327983, -802655152, 651522, 1456133524, -1395182473, 1888138},{2176, 67108864, 0, 738197504, -1135310447, -300696044, -156732242, 249561730, 43591074, 798693920, -688563309, 1294738},{-2147287040, 33554512, 16384, 1892679680, 986345857, -837323219, -957214503, -1350971892, 1904864076, 725373800, -282210738, 1080010},{4096, 67108864, 268435456, 590863944, 1277780849, -964067238, 1195110481, -813140903, -1592348405, -486469580, 168820760, 1070339},{4096, 48, 16384, 817487456, -61568335, 734883940, 2067592205, 336895183, 1506050, 425017344, -974826169, 968449},{0, 84410432, -1879035904, 1895120928, -782726983, 1586076578, -1252273196, 1281622038, -967815586, 1735074240, 98879068, 1301303},{0, 84444672, 16384, 819317856, -866454959, 755590690, 571838601, -796316208, -1663024113, -754847654, -2124609646, 384516},{327680, 64, 1879060480, 1898298720, -1859604039, 43296876, -610972524, 1498728709, 43341428, -513909532, 1441123983, 554697},{395392, 50331712, 20480, 301989888, -1151980927, 1993588260, -1905744242, 207681558, -121619951, 1992691864, -258406515, 495309},{0, 1729101824, 1342194328, 829926861, 1523354033, 1020037220, -1718941007, 412917392, 852136842, 1862658745, 1709377121, 823189},{0, 16777216, 344203648, 580653, -1224736768, 1023508, -439056616, 1192857756, -1868761964, 1855195465, 1824116615, 811736},{0, 16777217, 0, 21058560, 927351552, 1539629, -131694592, -1359182066, 2048439049, -1032220944, 127674064, 1466774},{2048, 83886112, 16384, 825743946, 1170509485, 1758275105, -1224016783, -1981191668, -1911784792, -211150619, 1251315292, 606150},{329856, 1572864, 268452608, 817537065, -381896551, 1502423720, -1956251297, -1879018425, -2700935, -152045676, 2006188054, 551591},{0, 48, 8192, 1107296256, 2043038386, 752539, -1369912828, -852200426, -841132375, 886380868, 423677389, 718549},{0, 83902512, 16640, 1644167168, 2084616305, 1023125, 1148800016, -591085296, 2026771104, -1506890386, 803013781, 1418968},{262144, 48, 402661376, 452297395, 1622184521, -2087823837, 861687209, 161248397, -2084094310, -1332066487, 208717709, 1495704},{327680, 101220400, 134234112, 1902739793, 1548261545, -1839975714, 1798148821, -1831234873, 722152191, 1184951023, -651613424, 1886098},{-2147287040, 64, 1296179200, 419155392, 1277991089, -716074156, 1861704901, 1641663575, 1464626012, -640874832, 1073741825, 1516119},{329728, 33554496, 12288, 521207808, 1789214809, -1534477083, -2020054384, -1803245306, 1213366062, -80538903, 1246536847, 1112743},{340418, 64, 268444032, 821330605, 1801246833, -693359450, -674487674, 1195716609, 801547944, -2063216551, -265509046, 1888983},{262336, 16777216, 8192, 617676800, -1690791559, -1760077146, -409685021, 104071186, -795250276, -1016112604, 218653523, 1258332},{65536, 0, 384, 2424832, 649163008, 1641250333, 452427841, -1069285040, 21448033, 1080253236, 1714795328, 1493663},{-2147483648, 83886097, 16384, 1898298688, -1857767311, -816831014, -1117071732, 806990864, -1273384030, -7147435, 227278872, 1667947},{201326592, 83886176, 1342193920, 1899477357, 1531221905, 1440055384, 553256724, -1327598512, 755320636, 989975569, -446693376, 1449714},{0, 87031872, 8576, 652279808, 1691500921, 704043, -665419776, 1164824204, 1809530454, -1771704265, 911855303, 1071047},{272576, 0, 0, -995393536, 810705267, -1810516453, -1902926362, 1195650498, 763709524, 1224000220, 1330118661, 1084564},{0, 69746720, 12288, 1689878528, 1279572137, 1901023272, 1756057288, -949181753, 1439033173, -631884837, -2022921332, 389013},{2048, 0, 16652, 310411264, 649212089, 1888386261, -553077211, 421871698, 1451416, -2126540088, -531926823, 606741},{2048, 64, 8576, 579895296, 900371065, 1540800043, -409635115, 1459099855, 416635506, 559961844, -1490457337, 825033},{327680, 16777216, 16384, 369098752, 683710137, -2037549863, 1070549688, 1214775296, -741372245, -1680929472, -851402096, 1451988},{0, 84443136, 16384, 355958784, -617572215, -1978745706, -1731440439, 7, 2035274122, 1185659046, 818776531, 466749},{0, 1048576, 0, 1199112192, -145383093, -237937260, -1588935872, 1327284502, -296164114, 1184148116, 1073741833, 214209},{137216, 67108880, 0, 805306368, 89252009, -669950483, -1568198659, -943962297, -661717306, -1351000843, -943962292, 1418438},{-2147155968, 1572928, 201351424, 1855567956, 1490585745, -1592445410, -476820172, 661159502, 2025859946, -406358616, 1779791576, 1295017},{327680, 48, 1210859776, 523618641, 1281145017, -1727184804, -491926828, -2147483620, 1498913370, 1228673860, -178177200, 1894253},{-2012872704, 68681808, 0, -1341466560, 744262235, -2087479777, -1969615755, 1832306447, 1712763562, 315960865, 1448444874, 926054},{-2147418112, 67108945, 256, 817889280, -421857967, 1561427478, -1892952619, -1278649017, 743034489, 1469240265, -1294124011, 1067980},{397312, 85459008, -1744830464, 817595041, 1277210177, 495932012, -1027099164, -1070739647, -1861457970, 1725643977, -653262836, 1435650},{65536, 50331648, 1744830464, 10518946, 1547268608, 563330463, -636203447, 18, 1195376640, -1297822136, 1148527058, 1240280},{264384, 100663296, 134238464, 1895128078, 1545900697, -1470746078, 734815922, 1293734272, -775824622, -418640044, -1291514091, 1895381},{201599040, 100663409, 33816576, -323240627, 2084100209, 1913988626, 309783186, -1266257343, -1634966738, 1670432545, 1494064780, 675735},{272384, 16777248, 0, -1317994176, 1278072971, 898604186, -1685381060, 63982480, 1024099844, 1579636256, -1073741808, 160843},{327680, 33554496, 24716, 512753664, 1540143193, -1991629988, 462895937, -661022073, 878250703, -885156911, -97024039, 834415},{137216, 0, 17048, 815380544, 1186763449, -99504048, 503607324, 22, 1560281088, 419075541, 962787367, 159590},{131072, 48, 4096, 1902215168, 2084171012, 1269285, -1022787584, 380655888, 182141804, -1897755475, 1289554637, 1487449},{0, 48, 256, 1769472, -866281472, 949786, 1210960184, -1966342139, 1316596, 1085033196, -1331417591, 1025794},{201326592, 69730401, 0, -1340801024, 541895019, 1523297251, -931869556, -1519418354, 1904689750, -564582548, 210787084, 1515637},{134490112, 96, 46137344, -1321138635, 1639240305, 92941849, 318632953, -448073908, -284553683, 1554893528, -1862755760, 1241442},{-2147024896, 70254673, 1879048320, 817605314, 2085923225, 1342992, -967355880, -156169387, 566709077, 1050163125, -1518765224, 970411},{-2147352576, 64, 12288, 818652224, -1227292591, -837583332, 648759853, 759169814, 51379096, -171520712, -597109668, 1511366},{65536, 69828608, 8576, 486211584, 1549044313, -37644762, -687271980, 414449686, -1974010996, 1995947219, -1318745083, 468594},{0, 67682304, 0, -986200032, -1495875483, 1678472722, 149833272, 13, -484663296, 852770126, 238144083, 855140},{6144, 64, 4352, -252706816, 1275517013, 25924714, -1563646408, -941075176, 1427123811, 939640808, -80190437, 1101433},{-2147287040, 83886144, 256, 1589138464, 1277466449, 1989421612, 511103012, 1743014223, 285619950, 178344213, 1687683085, 1356340},{-2013265920, 87081024, 0, -1321743936, 1759284569, -808834260, -1757690520, -1115252265, 855644111, 912489867, -1815030373, 710973},{6144, 67108880, 8192, 1890169920, 1732966405, -826167777, -411535775, -657894777, 1384615894, 1465489609, 501307856, 661350},{0, 48, 16384, 807043072, -190684495, 769556, -987332608, -802094382, 55927539, -1358326991, 1364797125, 353084},{0, 33554480, 1744846976, 825739723, 1279563857, -124368850, 5934988, 1496643802, 1494107040, 593397160, -51380210, 1896135},{0, 0, 16384, 1891272320, 1277542996, -1445815334, -703299136, 1355612053, 487207181, 1224200056, 30714369, 1085176},{0, 50331680, 16384, 13632832, 2067395840, 1012175975, 487522704, -1010531251, -2076168451, -86668036, -1584081508, 1661790},{196608, 17, 0, -1832889344, 96389739, 1498586223, 1250350789, -1190395890, 1837994724, 1820986277, -2002732472, 84614},{73400320, 64, 0, 792186880, 291015313, 59470699, 1478938817, -255650781, 102097, 1681723560, 277678723, 162060},{264320, 1572864, 0, 488636416, -1700229799, -1986610216, 1785866023, -930611192, -1902530094, 262056633, -1658025767, 1487246},{0, 16777248, 12288, 1887469568, -1420645267, 617331602, 1130186688, 1148724416, 2076430964, 1992757844, 1381268418, 220922},{393408, 84934768, -1207943168, -256293567, 1545924481, 1493710364, -1550144114, 1332740118, -719788152, -1757562324, -662105910, 792482},{-1730084864, 66, -1742077952, 821410135, 1817753745, -37123942, -1359065120, -328269777, 1904506491, 1146621788, -1891631095, 371802},{329728, 1572864, 16384, 1881899008, 472157817, 1267439125, 929839172, 122702733, -611891836, -1360807868, -1073741808, 1657580},{-2147483648, 67108897, 4096, -356483072, -64640843, -318079460, -241087304, 1859125266, -2016751953, 1259026913, -860042352, 608063},{0, 84410416, 17160, -1317418944, 1196988537, -808878046, -385168128, 434688089, 181946112, -1485658759, 1733495753, 1588935},{399360, 16777296, 16384, -243728384, 1094318251, -1529455981, 789572264, -1133754471, 1905864431, -560459976, 477120458, 1236645},{327680, 70303744, 256, 22526016, 281580544, -1688814377, -626452151, 1495531521, -1748297317, 332183478, -1186098023, 1497687},{0, 87032320, 17292, 1461757984, -782448231, 1703837228, -2053974339, -982253543, -956726933, 1990520135, -50702524, 1187630},{266432, 84410368, 0, -268435456, -1252747133, -1961781780, -2029178501, -2067418230, 1847116654, 118088897, 1502085139, 313753},{69632, 50331648, 16384, 19234816, 1509949440, 768720289, 1046753305, -805306362, 22090179, 855940161, -220123698, 1668816},{-2147483648, 83918865, 16384, 288358400, 1279046033, -217400740, -1046816592, 714634314, -1706672540, 598974494, -1966825578, 310954},{268288, 0, 256, 469762048, 725721481, -162047329, 1115596564, 1073741851, -91460438, 1688881812, -1125065834, 496254},{131072, 68681728, 4096, -771751936, 1817275027, -1403544021, -553450780, -2058605238, 1515020041, 576120140, 1254662672, 1301082},{0, 65, 384, 817890624, 1815466332, -958941665, -1334409315, 1706058629, 1670176727, 75045996, 798070170, 1468383},{274432, 85458976, 28672, -266829152, 1227132852, 1788304028, 1244526260, -902534523, 1817430775, 1326936189, -708837361, 189296},{69632, 96, 134234752, 1899486666, 1245100213, 424433700, -1906658780, 328204303, 34041634, 691703845, 866714258, 373449},{0, 67108864, 20616, 830049824, 740604017, 22434755, -1736014924, -1011600299, 1103494, 1580482580, 567766160, 1452714},{196608, 67125248, 8192, 426835968, 650418353, 2026797781, -945973104, -949111997, 901959800, 517320958, 433435474, 104196},{-2147483648, 35127362, 0, 662110208, 1355322985, -867459037, 351393917, 954790159, -897568044, -1564838223, -590872568, 1606023},{65536, 67108864, 12288, 87392256, -1674914436, 1813091776, -1031874568, 240222096, -451959609, -1492474540, 89418840, 254591},{333824, 33554448, 268451840, 1890288082, 1280095401, -1370076642, -409261656, 162044238, 1246411338, -343374692, -1964507112, 1877658},{-2013265920, 50331714, -2013265920, 750486017, 1195160217, -1844106668, -1401859508, -1480121132, -171617666, 2134675276, 153354244, 1041654},{0, 84983808, 16384, 504791040, -1690789751, 14129828, -314354815, 1073741846, -1932071613, 396553559, 2026704138, 301841},{0, 67108864, 1073750016, 816568931, 1277542817, 1775218202, 19321516, -760452652, -791722202, -1026829320, 1292659219, 372533},{-2147287040, 557122, 24576, 671088640, 1789439873, 1548467747, -942368915, -1225523187, -720032884, -746293173, 1558802382, 1416912},{-2147483648, 81, 1396719624, 750378607, 1547998609, 1329244, 361725952, -1387998201, -1886205021, 1356091193, -101313078, 1208011},{-2147352576, 67108944, 0, 294912, 1977284608, -2070588443, -355332844, 1728064921, -2065894644, -342569696, 117714325, 693381},{327744, 67108864, 8576, 1891696640, 1278636633, 722828829, 1257499322, 1, 96644096, 1268682849, -161413567, 676423},{327680, 50331712, 1128402944, 20294210, 1201969152, -905005714, 530276973, 1457637901, -293058675, 999850776, -2089488757, 1658722},{2048, 64, 0, 805306368, -176072599, -753433060, -1080528623, 38535190, -1994846259, -519743020, 38797330, 1055181},{0, 0, 16524, -1317421728, -1858561963, 51218468, 1361397696, 355467266, 1393505317, -58965967, 1691035017, 162380},{0, 102236240, 1124089856, 1890141473, 1815910585, -1470732132, 1692109496, 15, -845337088, -1614534888, 933276568, 560942},{393216, 69746688, -2147454708, 455597504, 1783933873, -1723701726, 1319262501, 1485570050, -1744165480, -1088063045, 1789547783, 1432236},{0, 17, 16384, -973078528, -332883797, 769448, -1056013164, 1690585412, 344959658, -1055915684, -1514924604, 366326},{-2147483648, 68157457, 0, 1890615296, 1753356293, 253203999, -1057958439, -1361776426, -37401042, 1180331732, -707195063, 707421},{201590912, 80, 0, 1533650976, 1246271657, -2075427944, -1168431214, 1738738692, 705123232, -1585756092, -1029701627, 1284185},{262144, 16777216, 8576, 705298432, -1531407719, 1909947116, -741925488, 14, -716760064, -1418945435, 1973536330, 1513224},{262144, 84444672, 0, 1895128512, -1943753623, 1750279682, -1359296888, 1183318032, 581937268, 2067444263, 56371077, 1059449},{-2147414016, 65, 20480, 1903689728, -329680775, 872490, 1849386356, 2021676936, 811363892, -1130654967, 1237135497, 1864571},{4096, 16, 0, 9437184, 447308544, 1993522593, -1885493932, -1968897465, 1092325, -253439760, -1863256761, 698626},{131072, 64, 140, 824180736, -698838199, 1900772244, 386812576, -1073741809, -330991975, -520730036, -282944816, 1606602},{196608, 16777281, 184549376, 10068566, -1224736768, 97369172, -97664928, 868774999, 781925093, 1458325272, -2141192187, 520750},{65536, 35127296, 0, 1890615296, -332286716, 1997520428, -1419357308, 141033481, -187118473, -1572179768, -1655929148, 715622},{0, 50331648, 0, -1004994560, 1471535108, 703891, 1948616980, -2108124864, 122642186, -1288335292, -1811601644, 1092872},{329920, 67141632, 268435456, -256287184, 1814607987, -116055485, -213682450, 3932188, 1586467279, 1728919759, -577502186, 1505748},{69824, 83886080, 2059681792, 1097455188, 1277474899, -732858864, 119993006, 114032660, 1829536877, 924748936, -773273456, 1089423},{327680, 65, 24576, 1891172352, -257548207, -1953483312, 1859240901, -1390399524, 1447443320, 160159924, 1073741827, 1020502},{262144, 17, 20864, 24183072, 120098048, 80712791, -1442737984, 1885340166, 998100, 1695285328, 539036118, 1016342},{262144, 17825792, 0, 821329920, 1347194033, 1519874917, -1751605724, -1073741823, -758797990, 1317353725, 1563253512, 1783897},{262144, 50331648, 8192, 652969536, -866871215, 875908, 391398992, 277636352, 163755884, -203613079, 260134041, 1491930},{-2147483648, 35127360, 0, 817413440, -534734671, 1068522, -988066588, -1497031866, 484128622, 506983001, -808923517, 152860},{-1945829376, 96, 16640, -1318474080, 1545902187, -1378724894, -1290268876, -1120504746, -1705448547, 387467992, 1869195089, 1886857},{2048, 102236160, 134234760, 1891317832, 1252298577, 1189158, -903536640, -903011062, 622428562, 1987869081, -1302623796, 444154},{-2147483648, 33554497, 0, 805306368, 1722442073, 1900969451, -1147564136, -1587738166, 1129876188, -1559556275, 1400737687, 90435},{339968, 33554432, 16384, 1711276032, -1341504647, -577730468, 1325296828, 18, 1778819072, -883044380, 249093514, 599756},{69632, 1572864, 0, -1692393472, -1138405477, -1693008342, -1035178179, -2025484668, -1684825869, 1594897321, 1073741825, 912581},{333824, 104333344, 16388, -1362057152, -331567015, -1365886400, -1628377272, -1865896314, -1609640084, 248246472, 1977571917, 434959},{-1946157056, 33554496, 0, 1879048192, 725227586, 1547235, 1281540096, -1212783911, 1657603898, -1565900068, -810969851, 1099514},{71680, 68157440, 0, 0, 1766154240, 1846771165, 2010523413, -1929551076, -200688336, 1406758236, -1891537334, 358613},{0, 118489155, 20480, 827837920, -1596920975, -250792430, -1949659416, 1868038150, -838673751, 1312193704, -820720103, 460526},{196608, 524288, 1073741824, 16827394, 1738952192, -2003330347, -1221719020, 38832279, 26271991, 177994952, -2145861229, 1238485},{262144, 84410368, 0, 1425375232, 1255713209, -37644772, -1560932112, 1410673820, 1397643779, -351330207, 1410334734, 13651},{399360, 117440592, 1342193792, 830058191, 1948637329, 1754302634, 447703736, 1788084240, -1956850964, -479819079, 2025875666, 152234},{327680, 16777281, 24576, -264601152, 1487179701, -989160304, 852921428, -1213676224, -891997460, -351610980, 183015874, 998102},{0, 50331665, 0, 12301312, 721420288, 687645, -845625328, 614569541, -2125186091, -632699436, 1151441168, 1469177},{0, 33554480, 16384, 605454336, 2066085233, -888512985, -1435693692, -1923297200, -711719224, -1901426096, -1968908144, 349037},{262144, 33554432, 20620, 1559962624, 1162385569, 739613402, -1762056120, -1899727804, 180460, 1401651200, -40137763, 374639},{0, 67665920, 0, 823186432, 959040841, 1489631, -711344128, 1372951313, 440849178, -959925781, -807822826, 1103116},{329728, 68157440, 12288, 771751936, -799491967, -485319594, 1188177773, -2015563960, -275150450, -1573864648, -588976382, 253530},{-2147221504, 16777249, 0, 671088640, -1539534447, -27944238, 520894144, 814844423, -1983898110, -1009115951, 1487142934, 1957324},{0, 0, 16384, -2037380672, 281729210, 1351834593, -1429076140, -833587899, 702592, 273727488, -2012687791, 496236},{0, 64, 0, 1176174592, 1882571330, -1865188699, -2063495000, -1965555696, -1869053194, 420008008, 152080519, 1147147},{393286, 118489088, -1438629248, -254027157, 1277751697, -51368424, 1449947574, 1197998085, 1515430007, -216210004, -1521404601, 1059498},{0, 18350080, -2013249536, 821406434, 1455980611, -900304279, -453408723, 1073741839, 1904750026, -2019069788, 195869265, 634506},{-2006712320, 0, 0, 0, -1136833024, 1020368416, -886467924, -1429527245, 1673113, -1062387712, 181681420, 435498},{327680, 33554528, 16388, 360241664, -64710567, -1999724310, 1939495317, -2143274937, 962121530, 926548036, -107023404, 552697},{272774, 32, 28676, 1455431744, 2083032505, -575325588, 371564662, 222863433, 435053, 1224097792, 822043469, 1209036},{196608, 0, 16384, 504725504, -783774055, 1490274, 192925872, 1121782862, 1451926614, -1157965488, 402715545, 16982},{-2147221504, 80, 0, 1879048192, 1224898571, 1196513432, 1185851644, -1605278835, -2078736628, 1490042965, 406865805, 1456272},{0, 67108864, 283385856, 525742, -1177253376, 1272007660, 828049424, 1383091165, 655289691, 1741902065, -1889763003, 1659859},{0, 67633152, -1342156800, -256131767, -1941402108, 546072704, 1230537297, -1786175339, 1699108180, 1391735524, 1894054400, 1075054},{65536, 83886080, -1274789620, 595184107, 1547262121, -1743508654, -1421800215, -1791649700, -1815022898, 791368365, -283693347, 1422062},{262144, 32, -1342156672, 1803139107, 1212462225, -1811261410, 1396480393, -734422522, -1709350001, -644262859, 1943615507, 1395502},{196608, 84934672, 17152, 1528889344, -1337682319, 685210858, 47579796, 1197998097, -981453271, 1532194012, 1817736978, 846373},{65536, 0, 0, 1476395008, -1185272491, -2108703524, -1172880120, 10, 93184, -1031845952, -2014020584, 330882},{65536, 48, 0, 10533920, 2069217792, 1313576483, 1465765645, 1212678156, 823634602, -347125687, -2008469238, 1433803},{0, 1124073536, -1171501052, 1894102345, 1549047977, 1058336, 2087800812, -817597352, -155099253, -688646020, 614615653, 91033},{-2147483648, 67108881, 1352814592, 1529167214, -1671907143, 1384960, 335544320, -1328966841, -112369811, -552743224, -1352331819, 973528},{196608, 16777217, 0, -451903488, 1548867692, 630631967, -1018309355, -183124926, -1135687036, -1091615183, 350299608, 981091},{196608, 32, 0, -268435456, -423018236, -942692842, -678817252, 1165281233, 2110891902, 892390149, 1393369616, 1680137},{-2147221504, 33554513, 4096, 1832365792, 1465166481, -1278711790, 785255929, -1380182586, 405475, -421799108, 1308367239, 1677006},{-1744830464, 33554498, -1476382720, -1552306496, 1454938236, 614484, 268435456, -1518691124, -1047937232, -1425502036, 1255981533, 1961734},{0, 68681745, 0, 360120320, 1152684721, 4955690, -1476016280, -529762491, 332469888, -488279840, -2147483636, 704000},{262144, 100663296, 20864, 458752, -1867881984, 1024730, -1979690416, 1096623368, 9479284, 453116284, -1348725248, 793368},{327744, 64, 0, -1331983744, 1279178909, 462564892, 1651995566, -1044321152, 1009173, -468072164, 248025552, 104470},{0, 83886112, 16768, 1131003552, 742498388, -61972963, -1467891648, -2145910765, -2113361279, 1805228188, -274726506, 429754},{0, 33554496, 140, 820366656, 471936353, -1202238289, -782004919, 1097864662, 1093230, -703194232, 1674819722, 1221419},{0, 68681728, -1342156800, -1322940798, 1280610234, 880674, -1265795072, 29627856, -1916701673, 372860260, 90707464, 1021688},{-2147151680, 64, 134217728, 1894493942, 1012048009, 84778533, -760270634, -1386650618, 821972, 1617281024, -1050647034, 857117},{0, 0, 8192, -2131066880, -1202642605, 1220130, 9280452, 18, -1136271360, -1268922903, 1376030149, 1573723},{0, 16777216, 0, -970227712, -1404502004, -796169454, -530234215, 29715536, -795412451, -412346775, -1050654250, 1021268},{327680, 524288, -1596833536, 828878506, 1279301745, 1858872858, 986859248, -2051014629, 1544365173, 936617816, 965056029, 372496},{137216, 16, 172244992, 829927125, -1462697855, -1861389084, 1264101640, -1995321195, 415549, 1819385096, 1497927887, 1492889},{331776, 68681744, 25472, 1663533056, 1792865905, 1988778016, 1456385372, -1983865913, 1316552, 254503360, -1567066363, 861804},{-2147483648, 68681728, 1207980800, 1865892962, -598176879, 22040, -841498624, -1473192755, -2095471805, 188595672, -36055031, 594678},{65536, 0, 0, 10518528, 962208256, 1397472797, -1759817535, 279713218, 1402331404, 1925957065, -717726585, 444445},{272384, 0, 8576, 470810624, 1515490129, -200332122, -1501372050, 1405172636, 721819745, 423068340, -125818042, 96791},{0, 67682304, -1140830200, 821803370, 721795242, 1829346851, -787904812, -755755568, 1069995327, -1025985289, 790240844, 436062},{262144, 16, 0, 103088128, -651022151, 1657502630, 1046676212, -1793764145, 407858927, -600173236, 353900618, 1045029},{-2147483648, 16777217, 0, 1140850688, 683865765, -1827955169, 25630684, 1930203145, -753952870, -564667695, 154522384, 1602989},{272576, 104333824, 88219648, -722088495, 2083862677, -2117327316, -1493502698, -2124677110, 1663572012, 1378758394, -1042016743, 1368705},{0, 83902496, 134234880, 485862130, 1415160649, 1901278506, -2000579972, -2026635248, -1379203289, 1124725518, 715702680, 293520},{-2013003776, 83, 24716, -1845493760, -1136297855, 1152532, -1106896536, -306310204, 1485992686, -1710811759, 1845467393, 530126},{262144, 87031808, 0, -1072037888, 473776810, 1758641709, 179014308, -1670555310, -951098197, -433753951, -596289198, 430184},{-2147483648, 16777281, 0, 425984, 1362923008, -1525959129, -1929718788, -1225261040, 1817523831, -354496355, 385656144, 1311024},{-2147483648, 50331648, 0, 87392256, -1807297164, 2009764846, -1736488920, -400010983, 98839, -1550873372, 1199623759, 522321},{-2147483648, 84934657, 16512, 1891336192, -1806520727, 1211052, 1093737376, 1790449174, -1170095346, 1511647965, -153800372, 809499},{0, 69747760, 25472, -756700448, 1414059673, 890529834, 1007113121, -1818230769, -2110796202, -1031837666, -256631737, 535120},{71680, 87146560, 0, 1459290720, 2084108457, -750083932, 1919839576, 336937217, 776489574, 310684331, 1322254355, 994546},{-2147483648, 50331712, 0, 17924096, 2066383360, 1925951013, -953822572, 1918745793, 1931001367, 1807555796, -2026779323, 1821993},{71680, 0, 0, 17825792, -111484416, 1812550182, -546410323, 349513025, 1297227976, 1661881473, -766246906, 1189153},{73531392, 64, -1207939072, 821803370, 1238935913, 1191248, -495610148, 1709072037, 1520158299, -2073109695, 1294494297, 1204119},{268288, 16, 21248, 1697972960, -1808232071, -942821216, 2138025193, 258765900, -939404532, -443234035, 1762971344, 1188746},{264192, 48, 0, 815846496, -1875549583, 525762072, 1053977025, 301280155, 1573345886, -1261040448, 5, 1226752},{6144, 0, 310788352, -1023693106, 1275181204, 1123864, -1567547392, 415029465, -809498228, -376697460, -399245094, 1094288},{0, 83886096, 134234112, 1899257430, -516114295, 798234, 469762048, -1967089463, -1408646507, -1362359976, 1891930629, 2679},{264192, 85458944, 8192, 1889533952, 683715425, 1003388123, 1390208537, 1412968658, 663237163, 199074144, 1077941760, 1934068},{65536, 67158097, 0, 580943872, -598701199, 1720687748, -1011295327, -1292257008, -1194407208, 505278919, 1449918473, 448954},{0, 87031873, -1136656384, -1338714047, -1136084838, 1620008476, -465938684, -1461703288, -1904207263, -1375444298, 1175191571, 1509729},{397312, 67108880, 268456320, 1890297544, 1522309273, 1434555934, 1248683397, -825666227, -317456660, -1977714720, 1632407643, 1805069},{0, 67108864, 4480, -995393536, 1280348076, -308917724, 96272440, 1222700434, 63627040, -541258024, -1461338936, 196433},{0, 68681728, 4096, -2068840448, 665360501, 1486331427, 41112949, -771895095, -792297369, 1470968317, 360448000, 1603537},{262208, 33554544, 1879069452, 729235155, 1428985961, 1926313252, -970153497, 388771675, 1422941, -832765228, 1746900738, 581408},{274500, 0, -1476373620, -248002112, 1280895673, -1376701422, 174420610, 1121981917, 282135800, -1852072683, -333534266, 302932},{-2147483648, 1048640, 0, 771751936, -1137405551, 1275392, -1458552832, -1343649128, -20594156, -1822870780, -1861717095, 1043850},{-2147352576, 100712514, 4096, 816918560, 406116465, 1355980319, -1171896300, -1562367862, 672992061, -1748537166, 135811353, 430614},{0, 35127296, 16388, -1342177280, -1709027573, 1473600166, -1604545223, -1787002858, -2145987245, -1629408492, -201171760, 170863},{4096, 67108864, 4480, 1891347136, -1673709414, 26365482, -1501384515, -2124677095, 965969960, 1933808553, 1949907649, 522833},{0, 69746800, 24844, -1355302816, 1438963345, 1989189674, 1215907748, 1406695053, 1079370560, 979151551, 857134549, 1391278},{65536, 67108864, 0, -1006632960, -173404747, -1999530468, -1575463660, 19, 1468566528, -2094656175, -1789831272, 118296},{0, 16, 0, 67108864, 1010717021, -1781088725, 549980468, 1230815314, 1316499, -1535144956, 497319837, 995106},{73859072, 67108947, 8192, -243780608, 1462546353, -627760556, 858126724, -1144013530, 429215471, -2045312612, -1049049471, 1219095},{201326592, 67108961, 268455936, 423048565, 1531492177, -1416345502, -418643492, 886447120, -1412231480, 840368604, 258743261, 603895},{131072, 16, 384, 23101440, -685135616, 949444126, -217426887, 1098913734, 186222171, 2080866673, 1881752448, 1502132},{0, 67108864, 4352, 16482976, -643480832, -762417770, -1049405756, 220749912, -2045404816, -1888188924, 1972930064, 1108890},{65536, 33554432, 16768, 403210240, -1479683479, -1488208470, 1789217632, 190952461, 677010, -493207552, -1434864571, 30302},{67108864, 50331712, -1795022848, 821415383, 1187289265, 664618, -1474412544, -121498098, 387290840, -286834204, 1319952346, 3815},{-2147483648, 1, 16520, 347718720, -599222599, 1599087936, 1706739753, -1587793663, 705173, -1333602828, 690109467, 677593},{0, 67108912, 20488, 806977536, 1456515673, 949586, 1880906632, 1104263297, 386078231, -413034496, -197165044, 492071},{71680, 67108864, 20488, 1903638208, 1549044825, 1867814438, -1883689267, 22816091, 148234281, -1492528999, -1147965477, 91968},{196608, 17825856, 0, 493453312, -125716391, -573211480, -1345501391, 285597123, 272984691, -426855927, -2147483640, 1510349},{-2147479552, 65, 0, -635764736, 744360819, 626234915, 1578493489, 1996039573, 418686, 1434550272, -615153253, 1497191},{4288, 69730304, 24704, 1860173824, 1799148185, 1016408674, 129825747, -1050935278, 1259971621, 869103953, 2040875783, 471694},{-2147418112, 66, 8576, 651538752, 1546043577, -796381660, 318283029, 1839258013, 1202028, -439271424, 720940620, 1408857},{333824, 17, 16384, 0, 2007617536, 1372689943, 1534259897, 700788871, 1675869, -1006632960, -1196600823, 862767},{201326592, 70254609, 21376, -335544320, -919811475, -691950042, -488845716, -1122525886, -959377509, -2104428076, 1852672476, 847505},{340032, 35127360, 0, 1453359104, 1012439225, -1727253369, -157534037, -644862319, 1406319196, -281005691, 1122512399, 1117079},{0, 1572880, 16640, 738197504, -1177249711, 1539612, -598769664, -1798811768, 1015180090, -433524555, 1939901954, 538152},{137216, 0, 16512, 17873984, -1682401280, 1837784292, 995619844, -1683392491, 875629, -630253696, -420365610, 1099356},{470089728, 33554499, 0, 1901702784, 1816478097, -1345445666, 438875473, 582359174, 1001276, 975883620, -1922772716, 1769515},{0, 538443808, 17048, 660684896, 1724427121, 412169684, 1688897984, -914313150, -1819015659, -1428819420, 1725594023, 1470394},{0, 17874944, 16384, 19945504, -597915648, 2139773842, -1134442984, -971210863, 394369261, 1398256934, -1312756267, 396824},{69632, 50331648, 16384, 1893743648, 1817598116, 274173479, 915793685, 9, -706913280, -1493757439, 1732059165, 591650},{262144, 83886176, -2147483648, 830048737, 1697419681, 1796388200, -637053227, -2040240626, 1716443655, 1061394136, 0, 896826},{-2080374784, 100663362, 0, 539394048, 1814867577, 701998, -563542296, -507314495, -19067105, 995727160, -709791673, 431214},{0, 16777248, 0, 1174405120, 1999970445, 1023149, -449376924, 1172624976, -742292722, -1288026652, 1403280912, 678156},{0, 85458944, 16384, -2059959904, 1421427034, -1936381396, 1693031548, -2000158706, -1403337495, -1821541739, -1701459962, 704230},{2176, 0, 12288, 1753219072, -1188385398, 747863452, 1454173026, -2147483638, -271647505, 70041968, -2124119992, 686614},{0, 1627389952, 17032, 1803103936, 1195151497, 1321556, -428228608, 1283724737, 663185624, 1987644804, -1364270866, 332417},{-2147483648, 84934721, 4096, 402653184, -425377703, 374311982, -1406188836, 815278357, 524860, 398145284, 386150291, 202262},{-2147483648, 35127296, 0, 805306368, 1010454892, 2094368287, -1870096423, 1732269064, -847130089, 327166097, -2059403241, 1218832},{2048, 0, 8192, 1882783744, 1705676442, 1527339, 1445537464, 310143874, 671891752, 147098689, -1941363316, 1507008},{264384, 83886112, 0, 1832205312, 1546016953, 1842261264, -1905050145, -2107820536, 1115965, 1665881260, 383867538, 1890838},{393216, 84410433, 0, 560565600, 1177062769, -1374710702, -2089964136, 561364108, -1131674008, -76549755, -922478777, 1020110},{262144, 16777248, 0, -637534208, 474560628, -950576509, -2044335676, -2147483623, -967203129, -1302428244, 96283604, 390239},{6144, 69730304, 0, -2059941536, 1549345210, 1325418012, 265381984, -964427759, -757545774, -1089701692, 1156868234, 550087},{-2147221504, 0, 12288, -1319106208, -333068205, -1277723558, -1214751943, 693755845, 604620608, -373044247, -1841299454, 1385150},{-2012858176, 67108944, 0, 1891183328, 1759021058, 932894, 730607214, 1843346573, 503711645, 1661518576, 62926600, 881420},{65536, 81, 1610629120, -252364512, 1547098269, 110116, -1829402312, 1894028377, 252257048, -116633347, -704835947, 1787501},{196608, 64, 8192, 1671168, -802646016, -2100593774, -876439111, -1741926700, 92058, -108542740, 1546502043, 1289937},{262144, 84410416, 8192, 344981504, 1464445793, 412333599, -160585336, 319652117, -2129165504, 779037357, 1096892552, 1814258},{262144, 524288, 8192, 423059008, -1672181159, -95326848, -1968320160, 1550915099, -972366432, 1714141521, 180199501, 1770082},{65536, 67108864, 384, -1321762816, 1278919354, 609325778, 129325081, 306446347, -1659764323, -764164295, -1151761970, 101926},{0, 68681760, 4096, -1433403392, -64106110, 1293732, 510017656, -2101859514, 730783503, 186396920, -1765474286, 1164141},{0, 69747760, 0, 595148864, 1431866233, 1900900394, 544327492, 1254126087, 540892777, 464875787, 1254922840, 1523037},{131072, 0, 0, 22023872, -1197129472, 1766825116, 979261876, 282956500, 1770415828, 2030947488, -2036807149, 971163},{196608, 0, 128, 1158676480, 1514760770, 492224039, 252461804, -1073741801, -205048786, 1694353176, -245035887, 431726},{6144, 33554448, -1119731712, 821803370, -1996343277, -2141808038, 1728999164, -1073741811, -1434065387, -1508468043, -1050663149, 1617449},{196608, 16777248, 0, 1476395008, -171845549, -846086742, -1703491391, -989544626, -1084570033, -1773157116, 1557921818, 944780},{0, 84459584, 402653184, 1902119351, -1406781348, 742930, 833978368, -513457388, 1531301615, 1043130375, -1822575147, 92507},{201588736, 17, -1342156800, 624405225, 1546948977, 1929620993, -91694424, 1737656580, 1933736664, 2041271204, 866989973, 582266},{262144, 35127376, 4096, 1891270656, 537524242, 1783846161, 120065168, -1797976812, 26042048, 103379153, 1284532951, 195273},{331968, 16777280, 0, 1526431744, 1345370289, 634280615, 1393653722, -968353707, 1686211199, -1575548932, -2139613102, 1425462},{-2147483648, 69747713, 0, 827343904, -1531317359, -1999913428, -1187374659, 763676803, -994934076, 647212042, -1066846830, 888891},{262144, 102236176, 20480, -1321874976, 1216419914, -828938084, -94678011, -1810618489, 387232350, -1622445036, 578672705, 98158},{264192, 32, 384, -805306368, -1135523436, -757678550, 1930983620, -1713791665, 68002307, 1694058264, -1214936504, 1118895},{0, 0, 8576, 1107296256, -180694387, 1661713958, 1555436129, -1044306423, 1661762499, 941343133, 966112329, 390748},{-2145189888, 66, 268443648, 1902140460, 473290833, 1268895, 2143847136, -1194929427, -1882198183, -468248155, 1098750402, 550460},{0, 50331648, 1342193664, 829938272, -1060805975, 1385002152, -468200747, -2122310384, 1385230687, 572298273, 1098727966, 678646},{262144, 16, 20480, -2080374784, -699090870, 1313569708, -879061672, -1050915256, 672188245, -209185452, 1360066882, 1868561},{0, 0, -2013265920, 1131907715, -1445637502, 1649128346, -1190346104, 1342726730, 684983479, 1889013972, -1047742591, 609010},{0, 50331664, 8192, 1098481664, -391550549, -1093691860, 1842814428, -933732516, 879354, -91912716, 1567407899, 1847239},{0, 67108864, 1218969600, 125403649, 658877267, 1467371, 492552192, -766164524, -2117649301, -1615493443, -689345008, 1314092},{6144, 83886145, -1207959552, 1899448747, 472430001, 730439745, 1655568088, 1993872849, 2038776736, -620655888, -2020857252, 716961},{-2147221504, 81, 268439808, -1341639633, -1707568828, -1114920282, -1163131067, 1006749574, -946709603, -126772223, -416956983, 1792897},{-2147483648, 33554432, 0, 1898010711, -1407111669, 1212915230, 1152406441, -1303117619, 587381519, -617851779, 22, 1191937},{-2147418112, 50331714, 0, 624404512, -597914767, 1330995372, 577978840, 1693739143, -2091136489, 1248383385, 1073741847, 478083},{-2147221504, 80, -1342177024, -1365656317, 1278523508, 1539483178, -960593148, -440626487, 1228557, 1885325612, -1410572351, 1686230},{0, 50331648, 17028, 821332640, 1540132209, 46628, -281001984, 1550666498, -716126763, 1728843933, 1892367761, 428623},{0, 69764704, -1879048192, -1321781897, -1068193103, -1673371578, -1934767400, -748680559, 656599832, 1119789726, -2147483630, 1425418},{-2006974464, 0, 16384, 805306368, 683003993, 676572703, -1448623376, 1694388339, 797415034, -240478916, 1156687876, 1298057},{0, 32, 16512, -1321959424, 1242104580, 1490274, 865917400, 1340967380, -1655240947, -1786687283, -132801268, 450070},{329728, 33554496, 0, -2046155744, 1179945835, 1737931732, 780740128, 108548056, 163901026, 2115621041, 279728149, 524343},{196608, 65, 128, 381714432, 682134953, -1898996323, -684026760, 599336084, -1885859059, 1696897473, 1954320128, 438985},{131072, 16, 16384, 1186570272, 1263048523, -1890944094, -362299276, -1661956266, 523878, 1650884968, 57153218, 402024},{262144, 80, 8576, 347834016, 1236918449, 1125279258, 1174672441, 1195683282, 1180409, 1621868544, 653045267, 245465},{268288, 83886112, 4096, -1317425728, 1149392981, -905108374, 1717495272, -2147483642, 1590957673, 2144887232, -861640256, 163421},{201326592, 64, 0, 807043072, -884587951, 1272558, -2009330680, -1214900388, 663132061, -1916270179, -1836793636, 717998},{460800, 69779488, 24576, 458752, 1430555392, 1461230, -426368204, 1340403717, -266583529, -1698026642, 29953862, 432664},{0, 524288, 8192, -960823296, -464409428, -804618734, 1552702685, 1557996437, 597197964, -1506907143, -872820647, 1871770},{274432, 80, 0, 1881440256, 566006705, -1169520553, -25134243, -611844082, -1413387339, 586432908, -609634092, 1099947},{67108864, 64, 134238984, 490188532, 1791538769, 1992917218, -1389869196, 895428497, 445380136, 1964396517, 1897343068, 1891980},{0, 0, 1879064832, 750332643, -1677068151, 550980, -2058102756, -1791131182, -1018005309, -1892871504, -1299944446, 1793719},{131072, 68681728, 0, 671481856, 984990073, 1381416471, 1914199332, 1159987229, 411708882, 937354828, 1096836295, 498730},{264192, 81, 268435840, 23713355, 1279045888, 93724, -2092834160, -369331118, -2037642645, -1810429844, 1791259778, 1502017},{-2147287040, 1048642, 1073741824, 528046625, 204254889, 1531532805, -80984608, -1296503664, 243369572, -1498467295, -790864254, 1343789},{0, 48, 8192, -1040187392, -701874084, 949804, -1670871756, -2107103224, 387711518, -263223128, -2105257086, 1826342},{65536, 0, 0, -2044035072, 934885444, 1389804245, 191761152, 34637323, -1093507920, 1805275748, 34637325, 632915},{272454, 100663296, -1476395008, -1665453022, -114155359, 435387026, -959257353, -981204968, 1505765465, 1732083756, -691447352, 11629},{272386, 96, -1144774272, 825608521, 1815654569, 657540506, 858137246, -689176554, -711354529, 14224769, -1403663146, 781872},{0, 17, 0, 3571712, 681709056, 1636457055, -1280452335, 1692946196, 1922828, -376367588, -1696493244, 193577},{262208, 33554480, 21248, 805306368, -1497052015, -2083561956, 716042638, 1256016661, 1217676189, 390158500, -398440297, 1108831},{262144, 18350080, 8192, 350997536, -1875864919, -1206490416, -423684328, -1954536124, 1649144177, -206868308, 4, 1737238},{-2147221504, 101711984, 20864, 1895148256, -532088679, 973942306, 655676333, 2042728390, 898285325, 797009721, 599525071, 1313693},{-2147413824, 66, 24576, 1845967904, 1791268497, 1720929824, 577217394, -1564644282, -1807354235, -1137948344, -2101046142, 783214},{262144, 87031824, 12288, -1342177280, -1337302357, 89619860, 1051575072, 1126170631, -942519526, 1535239921, -2032285733, 1343225},{340096, 50331712, 4096, -1687158784, 1764128849, 1582005144, -634667642, -1267173738, 1201068646, 1925864221, -618889533, 426590},{65536, 64, 20480, 1881440928, -1582526583, 2069020060, 998460744, -1743488172, -2124645674, -395211415, 1195213706, 468634},{0, 1157627904, 17156, 1691385856, 1881714297, -657744365, -923789472, -1073741823, -799579944, 840554472, 749103602, 4923},{333824, 68157440, 0, 393857504, -1867925335, 1871623256, 977054713, -1764187321, -1936554104, 935917996, -888360808, 1892719},{393216, 84410433, 12288, 1834024960, -801580927, -19825176, -1095270228, 729061381, 1904815856, -15732720, 459279045, 211725},{69632, 50331648, 402653184, 8469558, 616177664, 1229691567, -942804351, 1369994248, 1213577, -88096768, -747323445, 563336},{196608, 16777281, 0, 748781568, -531991207, 1838644754, 1594463993, -1559226789, 289450679, 2064635645, 1357381643, 1113361},{131072, 0, 17024, -959086592, -1805821804, 2060496994, 1919210960, 1461746385, 2061136976, -1541990624, 1736419074, 1289865},{0, 67108881, 0, 1509949440, -1478824379, -1957519854, -930690832, -1271361782, -1345146173, -1767291064, -927465460, 1321647},{0, 35127312, 268452480, 829935093, -802385783, -938560360, 883935285, -1963196413, -1886719345, 1310241504, 674875462, 328320},{0, 16777296, 1879064576, 514556579, 1548523081, -1403754332, 941462880, -2109123244, 1290051, -1767060960, -1035905534, 586554},{268288, 16777248, 20480, 716942016, 1221638289, -704481762, -146250068, 1185205704, 1905533850, -355020812, -1301779760, 93790},{0, 50331665, 16384, 1744830464, 992653962, -1034456233, -2000633812, 539803845, 704801327, -1418886488, 1814571656, 17960},{201326592, 65, 0, 1615936, 917394944, 949807, 56608532, 1994840075, 2046935846, -384971056, 1200424208, 809082},{0, 33554448, 268451840, 335988822, 1280087481, -1312064637, -170900247, 1528561666, -809132080, 798052925, 306040768, 790062},{0, 50331712, 0, 36339712, -1531589478, 767518, -726809432, -1273644839, -1191083051, -99017679, 472926934, 1616918},{393216, 65, 268455948, 787854358, 1520995985, 1329250, 1579500668, -1106910571, 1196571214, 1908808808, 2061680449, 1902481},{0, 1610612736, -1476377960, 515572290, -1675055463, 1327194, -1447591936, 404862867, -2113900204, 1100781973, -1584182411, 1806266},{69824, 64, 0, -1330610176, -1068910437, 735477290, -210654334, -1658301813, -1046710636, 676502852, 1073741853, 1918145},{272384, 18350080, 24576, 626623104, 1488306809, -1413380584, 525592304, -1652968488, 337411092, -1089132156, -893384893, 442885},{272384, 100712464, 8192, 1567671296, 1496617793, 1993297432, 668100456, -946309435, 1065533022, -1634426169, -946339833, 1502846},{6144, 33554448, 0, 1902166080, -1193424382, -1605198306, 588933864, -667417853, -918097195, 2114145432, -2147483620, 13513},{0, 557104, 16384, -250576896, 2082920453, 193633429, 807486748, -2122296571, -1537967588, -295765217, 1159728071, 1231780},{0, 87064576, 16768, -1021214720, 914503861, 621457, 145754000, 1200649931, 1078815643, -93788349, -1188521276, 342915},{-2013259776, 117440578, 24576, 1891347136, 1780797353, -1735290778, -1888081036, 938148237, 1904763425, -284360532, 99637963, 340741},{262144, 0, 128, 805306368, -1169866119, 1347591594, -615935096, -969406253, 327779, 1007206400, -225859578, 724847},{0, 0, 0, -1003028480, -63544907, 1544183314, 277087368, 1533053955, 1544044930, 632686784, -997389544, 1046038},{6144, 67108944, 4096, 1899407360, 1631631193, -1496542101, -2028280199, -931397614, -2017135692, 508533580, -1799533674, 564061},{0, 67667456, 1817726976, -243806766, 1524140570, 1901348896, 1159223188, -1874329600, 267486573, -1961789697, -2142957948, 541188},{-2147418112, 69730305, 0, 1160234432, 1546431163, 364924460, -1496870675, -1326639678, -216587696, -1302172552, 1333264400, 588999},{131072, 18350080, 0, -1845493760, 474052002, -191709651, -212479656, -893053560, -1588240212, 1051719420, -1976995884, 708268},{262336, 33554448, 0, 8421376, -80136960, 1788040676, 1799498494, -792392698, 25754218, 1057685532, 1353711619, 7437},{196608, 65, 20480, -2132443136, -121462454, -1269580380, 998689009, -1481001900, 1022500, 276531444, 410623244, 713305},{0, 67633152, 0, -1006632960, -145902963, -1706469872, -86506735, -1718016881, -976167914, -1495863508, 1380712460, 202122},{264320, 80, 268447744, 628734668, 1428994153, 1107381802, -1235620849, -1841494905, 1960318510, -1423030504, -1660337534, 797231},{262144, 0, 4096, -961970176, 339853995, -695054867, 59523472, -1718091761, -1974493959, 1392119149, -2121164144, 501661},{395456, 84934656, 16384, 1084278848, -329405620, 1204778534, -70223074, -951844533, -859540000, -886840191, 1341129224, 1893119},{0, 35127296, 16384, -2098495488, 380018866, 2052225761, 676070588, 124256278, 1893141580, 867771325, 1478756188, 1794900},{0, 67633200, 0, -1006632960, 618532491, 1049337365, 686163380, 98320029, 1579038331, -31086672, -944745781, 295617},{-2006974464, 0, 0, -258955168, 1790873714, 1545763, 1083739028, 969638459, -1148993708, -1610605719, 459914120, 759808},{-2012991488, 50331728, 180617216, 830046516, 1462276521, -1143819308, -1369113163, -1523943737, 503762, 1182719444, 1572453405, 496093},{0, 1124073488, 1207976600, 284539213, 1275771057, 55324161, 2060880624, -2144005283, 8473289, 648630581, 659467299, 572039},{-2147483648, 1, 17024, 347832320, 824479409, 16475, -1603043328, 566337607, 1942461055, -797325504, -1523287487, 1869443},{0, 524288, 230817792, 2802706, -780140544, 835615980, -1248667912, -1830551527, -917240544, -1711054031, 1376595596, 214473},{65536, 68157488, 20480, 815824896, -709738343, 1026984, 843628544, 121943813, -1937630451, -1415286704, -703837927, 1207048},{393280, 80, 1222656000, 1891183151, 1281150529, 1674881196, 779692810, -2126512128, 1262497300, 31539324, 504646469, 1499054},{0, 67108864, 0, 817528832, 550363985, 13715613, -1381283712, -997457724, -1459519414, 39789333, 448301142, 542121},{-2147090432, 69779456, 0, 452320256, 1629804625, -1491962792, -362376007, -125754300, 1573273417, -7243133, -2147483620, 426276},{329728, 100663344, 209993984, 360296136, 1243910057, 1838055458, 377763733, -788987500, 1114895, -503014532, -75644662, 306760},{0, 0, 16384, -2036760576, 1356505788, 1098939921, 582763636, 68681751, 1200388409, 1277973608, -876001655, 784020},{272388, 0, 4480, 819036160, 2083032665, 410164333, 2067460171, -1862992229, 625114, 1708773620, -1251693553, 1546756},{262208, 80, -2147483648, 830029506, 1448389225, 202083218, -1089081105, -674390078, -2079766015, -845162427, -1740373993, 438666},{-2147221376, 80, 0, 1654718464, 25270377, 2072943767, -216681118, -103695930, -1176731988, 475618461, -598881832, 1601989},{196608, 16777280, 134217728, 2859121, -1716481536, 1040874394, -1359543008, 419189254, 388878, 516293604, 1503411776, 1104600},{-2147483648, 65, 402653184, 322419063, -599162287, 2030592064, -1123776692, -1488684734, 1587835, -199163904, -946855678, 369268},{0, 0, 17028, 1827385056, -777371495, -137254766, -1659432612, 1095502479, 1625498, -670367744, 588647257, 48722},{0, 0, 8192, 1087733760, 1104560562, 1633113305, -2008786068, 313532114, 1214719, -1872674324, 71939840, 1321481},{262144, 48, 0, -266730976, 20220820, 1599520089, -1367947768, 0, 1598134116, 699811340, -668354984, 312442},{0, 1097792, -1335734272, 355949995, 1545899177, -619696860, -595915847, 492424453, -1258254378, 575159839, 196991808, 1215413},{474220544, 50331731, 134217728, -1695851032, 1420356697, -1614639615, -1035195147, 942108901, 2076754870, -891692872, -637502333, 502489},{-2147483648, 18350146, 134217728, 1443517474, 1473809081, 1091738706, -60140500, -343069686, 1795719092, -1293522032, 68419591, 439619},{0, 33554432, 4480, 0, -450441984, 1187741230, 221027612, -1659091248, 751346514, -760572627, -1341041974, 1932985},{-2147483648, 33554432, 16768, 481001472, 1414568081, -1990813089, -775497247, -415397567, -716726658, -696623775, -1579835811, 589787},{0, 67108864, -1476390912, -1317414321, 1275443202, -594834559, -2076966871, -2114175207, 1058092980, -4947460, -1761747754, 718747},{0, 50331680, -1824387072, 21047360, 901688832, 1180089901, -796392464, -724023728, 1057084075, 189646980, -881244198, 501513},{262144, 87064576, 1342177280, 389532097, 1222034361, -1702256614, 1202832505, 27, 1142173064, -155114701, -998663224, 84039},{196608, 16, -1476378624, 830069230, 289967449, 1329173, 257638824, 182721174, -1370466447, 1883969284, 1301321665, 1199665},{65536, 35127376, 16384, 1879310336, -1530875991, 181897964, 126390485, 337981637, 1116880488, -471763167, 1440025946, 1903527},{65536, 68157440, 12288, 829010976, 1487241297, -951100259, -1357983947, 265289732, 320568595, 1873360637, -1670002931, 1751929},{0, 16777216, 256, -1324318720, 933667698, 769445, 1342177280, -744997179, 1426672833, -2101214228, -334153338, 1517387},{0, 35127296, 17024, -2097086464, -1143553973, -623930284, 738204521, 10, 1944576, 2143365832, 1610987227, 1394562},{274624, 83902464, 28928, 659013664, -1140696975, -1139715264, -338517305, 367001603, 1922581948, 524724559, -1196592564, 339644},{-2147352576, 69828609, 0, -1375731712, 1700309889, 958570, 1983595552, -1555750127, -909051942, -1145659390, 1143284507, 826419},{0, 17, 16384, 16777216, -1404791040, 59478978, -1986061860, -117424499, -1713766532, 1192120497, 65799128, 1819343},{460928, 83, 16396, -248141120, 1817507985, 780676050, 911882707, 1675112064, 558668291, 352637673, -1134659244, 880519},{196608, 0, 16384, 716941920, -1866579279, -1387433944, 575216285, 450101253, 299019, -998505480, 130301831, 341930},{196608, 104349696, 17024, 1879411104, 2084083577, -1416454632, 1376322741, -983039993, 1457174614, -1757371654, -225686628, 1239840},{2048, 48, 16384, 786795040, 1255704977, -1236636896, 1939716137, -2067005167, 557929037, -1274999896, -1951915699, 299740},{327744, 68157440, 12288, 10507328, 1170249472, 613389420, 1059631795, 130579398, 807096347, -1240911288, -1023378300, 281409},{262144, 571998320, 402674432, 1559615575, 2025100113, 799332, 257540096, -855806528, 1841598347, 733375741, 1997699832, 558724},{0, 16777216, 16652, 822116352, 397973321, 760981, 2013265920, -2072229756, -1193450708, 1387251956, -38385509, 1198779},{0, 67141632, 4096, -1342177280, 470407188, 533703875, 1702711320, 1473536597, 26553686, 1249684895, -2113929216, 1704546},{274432, 83886080, 128, 1698004992, -516045919, 36378, 449291552, 1486618628, 412964295, 2072626468, 2023495812, 1323627},{65536, 1048576, 16384, -1330928016, -238512883, -909040382, 934576177, -1073741807, 878286062, 783268280, 253292885, 1402826},{0, 67, 20608, 1089845952, -1408870389, 1083522, -469762048, -257147325, 525387265, 2024670184, 1892949835, 439198},{-2147090432, 83886144, 12288, 1397784576, 4113081, 629901981, -1172225440, -1179113977, 379297716, -1639464423, -781647844, 1953313},{196608, 68157440, 20480, 485851136, -791890791, 1795854360, -1487158504, 89653268, 64423064, -414326004, 1185961347, 255595},{0, 68206592, 4096, 818971200, 2069139017, 1162501095, 632757324, -990356332, 828076484, 323238691, -2063836030, 294469},{137216, 67108864, 20480, 1898283008, 1354364420, -44608927, 383332600, -973602813, 714336, -1547223040, -972005489, 1682184},{201654272, 65, 25472, 313085280, 1791284921, 2123659360, 386753517, 1999011142, 126887, -1585741308, 1742479443, 1798911},{327680, 68681728, 24576, 1679196160, 2084866649, 1918257281, -156743824, -2147109179, 1127084, 259630968, -2027392442, 312951},{-1945829376, 67108960, 0, 820369504, 1429510329, 1862361254, -1301035224, -1544576953, 277328710, -490593227, 1144328325, 1681852},{196608, 0, 4352, 18926656, 1732681728, 1530515, -1366982656, -585087203, -2054382292, 541531672, -221126243, 1974},{131072, 0, 16384, 479264768, 1473053009, 1222032919, -1038237212, -2147483621, 1225259148, 721027788, 1207733463, 268046},{272518, 100663312, 0, 1566031872, 1496617817, 888222360, 1876026334, 1390994564, 1115895617, -825630152, -1940389870, 145636},{266432, 104349696, -1207939072, 816328239, -799500175, -543873518, -744850957, 124547329, 1229440122, 1115319698, -945786809, 120799},{-1744830464, 50331714, 0, 1608256, 1463588864, -2029431600, -631843968, -151041661, 696513055, 441160857, 312551058, 554119},{272454, 100663296, 8192, 16792608, 685541632, -1384948203, 1715414163, 4, 482462720, -2038662512, 1522008392, 1745485},{131072, 64, 4096, 22033440, -1808084224, -2146477394, -1167915792, -507960166, 84566, -192937984, -1044820476, 310050},{262144, 85458976, 0, 548470784, 1546172537, 600156, -1416887844, 1073741825, -1207954936, -1296388859, 30673028, 904120},{0, 16777280, -1744818176, 1892375970, -1408870307, 599554, -67108864, -1453304500, -658079108, 43388304, -984302461, 1320519},{134217728, 16777280, 0, 515407872, 1544143689, 538334723, -803878719, -308407167, 542867309, 36587717, -1050924966, 1402919},{-2147221504, 33554512, 0, 1882488832, 1495831385, -2075155558, 1396964693, -129386875, 441011888, -1820075868, 1533549131, 1885578},{4096, 50331648, 4096, 821803720, 1277850957, 587965979, 1736270885, 1077166677, 1142536244, 1271534132, 17, 1131076},{0, 16777280, 0, 1190513984, -653934070, 1458222, -1517268392, -1644848679, 634931167, -405224467, 25, 256063},{0, 64, 20492, 1578644576, 1532792393, 1151142, -792772608, 35397889, -1085132163, 405160588, -1130225200, 272113},{69632, 0, 268452480, 1895505987, 1422438761, 1066642716, 2050908544, -2147483637, 1447999, -697613548, -150454128, 15934},{329728, 1097792, 0, -447237088, -867919780, 265201152, 1311126548, 1073741840, -1220045296, 1780589087, -2105795247, 1321028},{0, 67108912, 20480, 818937856, 1631885145, 1091207261, 633471544, 1110966300, 719396, -98286572, 1895631299, 46699},{329856, 0, 16768, 1894809600, 1616687433, -1014342127, -1816708017, 1073741824, -1742985042, -463598860, -1112252795, 1216069},{339968, 67633200, 8192, 753631232, 1781830033, 2005555242, 733375176, 1293428376, -679085399, 387196712, -2116802494, 398039},{-2147483648, 1048641, 4096, 805306368, -708798639, 1145752, -2011364892, 577241092, 1201361791, 1870406796, -1697637036, 516013},{0, 16777216, 0, 1155554336, -1406775372, -771008986, -315832791, 404488214, 549585920, 2053276168, 404750343, 469504},{0, 18350144, 8192, -771751936, 1548783187, 1465893, -1675821056, -253424574, 801409650, 172194460, 446169105, 1706526},{-2013265920, 50331744, -1379777920, 816399648, 1530957433, -2108410342, 1080279505, 611476486, -2108346414, 439141013, -1110696610, 131682},{131072, 69730304, 12288, 805601280, 816361081, 605335077, -367050196, 1, 973225984, -1974307783, -2110700607, 184863},{262144, 16777217, 0, -243826688, -1135692686, -1844529638, 1261982364, -1176916709, -1840362942, 981949136, 2, 1215488},{0, 67108880, 256, 771751936, 1155041921, 948970, 1476395008, -671853563, -2071485569, -162150324, -138115903, 465887},{0, 67108896, 20608, 654029856, -2142717839, 1560456748, -1067678468, -825229311, 1350188, 2120008956, 1657859396, 1687175},{201392128, 64, 8192, 805306368, 1187672401, 752552, -1814490924, -1580213862, -1526375859, 1695369992, 281325788, 1753630},{-2147477504, 80, 16384, 1891183136, 1454937785, 1136763050, 793715776, 764203090, 1841678896, 1411553001, -1784676347, 327202},{266240, 50331664, 0, 294912, -172665344, 265643228, 1993997741, 1340927388, -304479473, -2111323812, -978583525, 973915},{327680, 68681744, 0, 438697984, 811382345, 1004453, -297156116, 1508216835, 516514692, 113031240, -2069870142, 1923532},{-2147418112, 66, 0, 808880576, 935745457, 130635281, -347897716, -514030142, 134219702, 1027342476, -2124380716, 166466},{0, 32, 16384, -949518336, -1875238508, 1399440, -864043008, -997179000, 2144989758, -1516681012, 1142685721, 1820233},{264192, 1097808, 134217728, 661077737, 738285657, -682267903, 1514305732, -637479096, -796090840, 1260610626, -756440957, 1321278},{0, 102236192, 17024, 715752992, 1689826425, 813092, 337446112, 81639427, -1205994645, -1814481135, -469915132, 523916},{-2147155968, 33554449, 16384, -1341620224, 1705023562, 1277413, -363980860, -445546478, -2146340319, -567818895, 398983175, 1317454},{131072, 85459008, 0, 1899472960, 1355331161, 952361, -97104784, -613664829, -624441590, -1774145284, -1073741820, 1844442},{262144, 84459552, 0, 425984, 1161597696, 926892, 1845493760, 1208241989, -1585379746, -1153260462, 1157136580, 716928},{196608, 32, 16384, 637534208, 270680489, 646558685, 984239388, -2130095166, 149009, 0, -1055566848, 5804},{340096, 68681728, 0, 1880653824, 1498188377, 646477842, 52739130, -945522168, 847456295, -136611120, 95967940, 298105},{0, 1048576, 16384, 817465056, 1814598033, 633029, -732838800, 1148190743, 1376306464, -1965579772, -1844961150, 35468},{0, 64, 0, 102467840, -1723977615, -1899340250, -441024092, 1542717456, 294426, -1716074256, 86884314, 126506},{-2147418112, 69730305, 24576, -2056700256, 1422166619, 1989424672, 723666816, -489841274, -950603232, 109866104, 1283269074, 1403492},{196608, 67108944, 1207959552, 1458275968, 1455724177, -2108927830, -12345976, -1002692734, 1796901, -1505867736, 1, 1294630},{266240, 83886128, 0, 814810688, -1137055079, -1240023510, -1167836711, -1994653671, -1241343297, -1574325331, 200839644, 250171},{196608, 70254592, 20616, 1894501408, 1154013363, 2039824418, 1114326352, -2019788478, -792179329, 1581166128, -1573753966, 256543},{262144, 83886128, -1342173184, 595052898, 1543583825, -1363118576, -138098396, -920342837, -1592077745, 1732901856, -2050190782, 1221566},{0, 67125296, 0, -2063597568, 961842061, 949807, 0, 1258832192, 1121437453, -1232804514, -2076687546, 677953},{0, 67108912, 0, 807961920, -1153922647, 1277412, 181984108, -690207805, -1224354091, 1984431229, -2071986149, 1418302},{0, 67108864, 0, 807960576, 1152158329, 1196134, -585477020, -1898101170, 1440586523, 376623544, -983826428, 470327},{0, 50331648, 0, 1157300224, 281608346, 306869099, 1225068621, 1564070616, 1242584338, 735419596, -2147483646, 1005011},{331776, 67125296, 134217728, 586502194, 1188337777, -900510320, 2064645289, -1649554809, 387825541, 710667998, 7, 0},{0, 32, 384, -2098180032, -1948856213, 654941346, -1848688227, 1207815940, 1592218, -130837904, 586169564, 304031},{-1945698304, 80, 17152, 1879048192, -247162735, 1096007042, 596006065, -1470135651, -2038431180, 1053873193, 942230356, 1581869},{131072, 64, -1595670528, 829882913, 908630105, 1250801195, -836304432, 1114947528, 123756, -1203060736, 1155579844, 202789},{262144, 48, 4096, 505872384, -601320535, -2024359232, 651650416, 153392728, 1306250, 0, -1993828736, 1706631},{-2147483648, 1, 0, 81513824, -1870514093, 534099088, -393130204, 1642107265, 538383274, 1955696372, -1893203956, 896030},{0, 69730305, 4096, 392167424, 1548257945, 1518178, 743391232, 587526346, 902132608, 646408944, 9, 1559040},{-2147352576, 17, 0, 821788672, 1504072771, 1471131, 644122928, -518780260, -1823408585, -1364556216, 181141517, 861231},{196608, 16, 17024, 808091648, 1547483289, -1064394716, 237524300, -2059403256, -1060633016, -1384458932, 632925509, 972333},{268288, 16, 0, -984138048, 1277802644, 411125266, -502210188, -765452479, 883222, -835551232, 1073741834, 1205279},{-2013265920, 64, 0, -1318633760, -869391508, 175636, 1409286144, 1663704836, 349818, -1172110804, 469350597, 1797151},{272384, 50331648, 136, 1899274816, 1280882873, 1146170906, 2115369432, 8421442, -2142472125, 172164160, -1307965374, 1563276},{266240, 0, 0, 806617088, -1313305183, 1103701204, -300260292, -2017161407, 2088787068, -1639857268, -2147483622, 232591},{262144, 83886080, -2147458944, 825724610, 1438177465, -1056099228, -1904712984, -1071644224, 189633, -2101379040, -1564463872, 273186},{-2147483648, 536870945, 17024, 781811712, 123254889, 1021009, -59686448, 603833603, 629426137, -1178267660, 876553766, 269887},{0, 17, 16384, 808878080, 2084664913, 1917754531, -1641561631, 1999110164, 1719918410, 674398853, -2115232119, 168488},{73400320, 64, 20736, 650182656, 1548268649, 1993324061, 154961172, -1482719253, 1998291683, 1011975436, -1428077612, 261739},{2048, 0, 16652, 817922048, 1698343273, -300450665, -292391368, 1327780106, 63209540, 609272708, -1134858673, 164798},{0, 0, 4364, -2147483648, -424760158, 1031724, 1498677248, 360448003, 470360, 1095991296, -1540147179, 268867},{196608, 524288, 16384, -2063580064, -600640931, 949798, 1107296256, -2147483644, 1923317, -2099692336, 1331443524, 387845},{-2147483648, 16777297, 16640, 1660977152, 1546687891, 24104, 1713183220, -1524629484, 1329753883, 799087116, -1129557433, 1393434},{65536, 69730304, 0, 807698432, 470112345, 1077443, 640303568, -1997537263, 1915434, 1850270520, 150253506, 1898522},{262144, 84934656, 4480, 1889533952, 1438248369, 1308732964, 1942660677, 127664132, -2105129650, 595976933, 567572933, 217051},{0, 69779553, 0, 806617088, -1672967591, 1422428, 975437824, -1473749053, 650289711, -217144354, -1037017144, 160898},{0, 84459520, 16384, 19237344, 1262786304, 939552, 613531648, 1544405129, -1844938314, -757598102, 2047456834, 411467},{69824, 67108944, 0, 1899331584, 1154791505, -1853327324, 460416226, -2104140989, 696384239, 706645392, -1030661176, 889046},{264192, 100663376, 384, 620759680, 1470927257, 898250282, 1653222020, 395334235, 597679, -567884540, -1526967655, 555670},{-1946157056, 64, 0, 1881594912, -1482609148, 761380, -330543656, -1380798646, -578269551, -861156844, -2067475830, 993868},{262144, 85458960, 0, 1891205120, -784770927, 542224430, -27572027, 450217156, 1224936375, -823056968, -1844969467, 1799308},{262208, 48, 0, 1140850688, -1529752733, 382688682, -690511110, 1210843152, 574691930, 485593641, 1378386703, 1163501},{6144, 67108864, 0, 816555712, 1145692825, -821122974, 796605685, -1807946109, 748178895, 1938086577, 250085403, 1749315},{331968, 67108960, 4096, 817431264, 1546988681, 134904720, -568876658, 487706766, 1548672604, 1607687472, 1170592005, 209875},{327680, 68206592, 4096, 1563754496, 2025107521, -2000061267, 1249679945, 1080108888, 127904, -1574755238, 1073741828, 1834791},{0, 50331649, 0, 1802240, 396741888, -305423211, 550997780, 583019008, 683946564, 1244564860, 30670852, 862449},{272838, 17825792, 24576, 659554304, 744159305, 1106324995, 1939499006, -2069043182, 1200081445, -1908114808, 78752003, 300608},{0, 64, 4096, -970534912, 2069171860, 1005075, 1476395008, 579174417, 1321474, -378366212, -1854605759, 795516},{-1946025984, 67108944, 0, 805872704, 1162655833, 1972272676, -27342824, 2085779203, 786175, -1357901588, -2011397756, 388190},{262144, 48, 0, 807994752, -534472551, 1343511194, 1935937252, 1186463749, -1044171901, -464565216, 1186725910, 795011},{0, 67665920, 12288, 622592, -1256114944, 965484, 1073741824, 154428612, 1146334548, 38908990, 154690754, 724795},{0, 16777248, 16384, 1897179712, 1368053947, 555929, 603979776, 202200332, 993238, 385240104, -334408443, 326202},{262144, 83886128, 4096, 653920800, -1672959399, 524322304, 1262924388, 1386226694, 634749738, 925254137, 9, 222720},{268288, 83886080, 4096, 1561329664, 1428984737, -1895733084, 1312269112, -2124677099, 172470, 265691536, -2118533428, 1124906},{0, 1048640, 20620, 805306368, 1196028313, -1676857938, 74684873, 1360367825, -465439186, 1335960272, 2046715011, 1205842},{0, 68681728, 0, 1881899008, 5849436, 634295827, -125659539, 184379080, -1886698316, 1857036916, -765460453, 576870},{69632, 64, 21248, 816873472, 1497743481, 462921129, 1196305397, 226492422, -980941095, 1706495024, -383663909, 1695431},{0, 35127296, -1476378624, 816546241, 1246040209, -1680650850, -1797714179, 1168136066, -1311208295, 1243837884, 186407362, 588700},{0, 64, 0, 806685056, -776283975, 1376943190, -263207664, -1433120694, 785312, 1486880768, 190337611, 332881},{0, 68206592, 1879048192, -1340451776, 400427293, -1303667563, 741457928, -1070858099, 1284364460, -1160171734, -1960271994, 205824},{196608, 67108880, 0, 1153138688, -1806548835, -1387631828, -1817371791, 95989975, 222125, 709379292, -996888375, 296013},{0, 32, 4096, 15765024, -1688844155, 1530534, 418217984, -2147483633, 718626, -872415232, 1369992337, 314137},{-2147483648, 66, -1342164992, -2060090815, 1195677114, 76030802, -1383804408, 1949901011, 75792964, 206193824, -2069625646, 1856463},{196608, 64, 4096, 1158676480, 1278310565, 599572, -1503896416, 1554895045, 470995, 735117312, 480630802, 1165259},{0, 50331713, 0, 1365056, -424488043, 1538772, 1890369956, -529428480, 1070980, -1281015808, -894952806, 233644},{0, 17825792, 16384, 823219232, -1531551655, 1226276, 25317760, -827557553, 988200, -942441812, -1892155387, 1879832},{-2147483648, 67108881, 0, -994377728, 604412012, 611651, 106939564, 1686658202, 233255, -94365044, 387711004, 1533302},{-2147483648, 33554498, 12288, 1879605248, 1087010933, 1462881, -1610612736, -1343974968, 499586, 2132167000, 194248717, 182970},{-2147483648, 65, 8192, 807075840, 539387985, 1385309, 1946157056, 695039831, -1387921495, 1079953436, -1995087550, 951959},{-2147483648, 33554496, 20864, -268435456, 1277725044, 1523421224, -446036695, -1407093866, 1938324338, -632120839, -536870889, 600960},{272384, 0, 4096, 1881585696, 1279871353, 2048089368, -359552716, -949454783, 2017961081, 40159100, 175678865, 532088},{131072, 1572864, 16384, 824180736, 1354012273, 2119154921, 717277392, -1073741809, -1941213066, 575714640, 1259372172, 338609},{0, 0, 4096, 1614187200, -1715840836, 679454, 1543503872, 308543489, 1338903, 2082013184, -2114453503, 1340953},{0, 1572864, 17024, 1881605792, -64362111, 1542892, 1559304004, 1445986305, 420414836, 1187160744, -1358692335, 1182348},{0, 32, 17036, 805897536, 1278646413, 632345, 1075746560, -1761607679, 1498588719, 1076790001, 575082631, 537111},{0, 50331712, 8192, 1507328, 1277726720, 1152426, -509584968, 667713031, 977433, -226698744, 189042587, 212839},{0, 48, 16384, 807829504, 1487765921, 1211805, -900380448, 1128290649, 1510884866, -1878899904, 1222639629, 34446},{262208, 0, 12288, -997195776, 1229755474, 487961498, -882448134, 7, 367616, -1541013504, -912523240, 721496},{272384, 16, 8576, 1678114816, 1471459697, -1730784665, -368956764, 1263271938, 1838752, 337903616, -353107963, 800539},{0, 16777264, 17032, -1342177280, -868812790, -7321596, 537237988, 1341420611, -1878053986, 513785869, 969015499, 155200},{0, 1610612736, 17028, -255819776, 1543649429, 478851226, -2073307083, 97255428, 479697273, 1517017145, -451522389, 166430},{71680, 67108864, 0, 1890629664, -78470653, 2098372066, 182302065, -1073741824, 675803262, 2001961608, 41974023, 731988},{131072, 524352, 20864, 1866465280, 1524141689, 1431409690, -744712200, -2069625638, -1856489667, -2041711555, -1307468732, 442285},{-2147151872, 68681728, 0, 1879048192, -1487292230, 1884380190, 1126022416, -243415339, -648964326, 1190261121, 1145834308, 1879513},{0, 16777281, 0, 10569779, -88464640, 1347862038, -1930260736, -529206653, 1925920, -1498625140, -989331452, 20139},{0, 50331680, 0, 56688640, 936046082, -1198891501, -1353835635, 1535901724, 1905396, -2098559116, 1073741853, 989464},{0, 33554480, 16384, 816545792, -1873657487, 1291610, -1796830984, 100437906, 1730422, -1826240472, -1073741821, 587484},{71680, 0, 16384, -2071953408, 273979499, 160611731, 397078897, -1047258865, 612583, 1879048192, 1, 412160},{-2147418112, 81, 17152, -1318486016, -601499479, 1151144, -1902720744, -498539366, 161649, 56727220, -173015034, 1204866},{65536, 67108944, 8192, 805306368, 1883276169, 1270957, -1424015360, -1846018040, 1795666, 593187320, -1765450871, 762734},{-2147155968, 67108961, 0, -1340538880, -598951822, 1989521536, -1820891960, 1692477197, 659930797, -1703426847, -947312830, 500812},{196608, 0, 16384, -265781248, -1602111486, 961682, -97417148, 41190681, 1522353, -239205608, 8, 337541},{0, 67108881, 20480, 607397920, 1152841841, 760812, 2135774440, -231997430, 493175, -886914664, -1049624572, 709454},{327680, 18350144, 24576, -1342177280, 717587049, 636125, -1148839896, -2147483643, 724835, -625509712, -1237744184, 1799806},{0, 17875008, 0, -2147483648, 1280870770, 861354, -268435456, 1171259394, 278014580, -2112265865, -1073741823, 166233},{327680, 16777281, 0, 1879048192, 1786919025, 444618263, 1333028812, 2077080728, -1285752080, 372874189, -1013327985, 1706397},{327680, 50331712, 0, 1879048192, -2134329342, 365922472, -948953044, -2147483643, -1214433609, 1183728456, 1119923713, 10292},{-2147352576, 17, 16384, -614432768, 958472277, 753181, -497427788, 1650497991, 1254608564, -1867392328, -1073741819, 109093},{-2147483648, 67633185, 0, 818946112, 1815803985, 1502567507, -378464511, 575184903, 1929389620, -1839582972, -2014807806, 583349},{0, 48, 16512, -603979776, -1858701133, 1400868, 1879048192, 1564070746, 728976, 967268480, -268894371, 308124},{131072, 0, 0, -971440128, 2057925708, 949805, 1717327000, -746061813, -397507477, -155035760, -1801715702, 796035},{264384, 83886080, 8192, 1879048192, 959012876, 1410626393, -274830537, -965738491, 165013, 525814068, 8, 206568},{196608, 64, 0, 539264544, 1186635897, 1479312, -883632792, 1073741841, 795331, 223772672, -1787297780, 1690944},{0, 50331712, 20480, 806879232, -333137775, 899234, 341884928, 638320647, 1321619071, -674561499, 308568279, 604952},{2048, 65, 20480, 1820360704, -869615507, 1539460642, 60596308, -355729384, -841657533, -1201844876, -2049910845, 791099},{262144, 84410368, 12288, -1328447488, 1094236282, 1203539, 1714012784, 1114374162, -1190899956, -69635707, 57941313, 1881017},{0, 64, 8576, 1638400, 1990642688, 948949, 704643072, 225252047, 174968, 1695731636, 848897548, 234169},{-2147483648, 33, 16384, -1332724736, -1137041068, -950641110, -1902797471, -1118447525, 1369835, -2050031616, 1353749149, 192025},{0, 33554480, 16384, -1040187392, -867919790, 881892, 1345388544, 1437954194, 382627691, -747597132, 1981622989, 1471350},{196608, 64, 4096, -1006338048, 2063947946, 814309, 2132777668, -624689138, 889709, -1515634688, 21, 1144668},{0, 16, 256, -2046820352, 1194677132, 1408535, 1957861864, -949209518, 1541751, -845211372, -349396476, 621284},{131072, 67633152, 0, 760217600, 1275667345, 1140250, 1001193472, -2102885161, 1305606705, 393128016, 5, 0},{0, 83886128, 16512, 826290208, -1253686631, 1471338, 747408136, -1758950190, -1375411687, 254240972, -148281600, 3660},{262144, 48, 8192, 805306368, 809277609, 1151069, -2021336416, 373402116, 1827718, -1476395008, -2147483644, 726602},{0, 0, 4352, 20975136, 1504276992, 1474077, 143163392, -929749167, 1191893, -1725480960, -278122686, 1366862},{201326592, 83, 16384, 1811939328, 1350714009, 600867, -863909132, -88928485, -1706777084, -520729880, -1325366950, 1184628},{262144, 0, 8576, 825655296, -1607630455, 1224232, 317882368, -1838153699, 724020, -1677721600, -1586419246, 383857},{0, 1097744, 16384, 826310656, -1135760799, 949674, 1615937536, -880017406, -1705259343, 2074125210, 93606109, 330330},{-2147483648, 50331648, 16384, -2080374784, 1275205770, 617321258, 74028041, -426164086, -1249150412, -897673460, -963117054, 990050},{262144, 50331648, 0, 807010304, -1606032751, 1595235858, -70024540, 99352584, 387314783, -1157654719, 274472282, 1523991},{0, 0, 0, 103186432, -1430707843, 1293732, 1101250560, 1073741850, 1116866, -1726558164, -990046502, 1545561},{268288, 16, 0, 491817376, -1138405564, -414083604, 1268705244, 2, 1915392, 1994866688, -1073741798, 517354},{262144, 16777264, 0, 823164928, -1856678815, 63664976, 724239116, 51118085, 625903445, 660050957, -759879476, 1351488},{196608, 33554496, 20608, 1879048192, 1549572169, 618015258, 1920795476, 1741709382, 1619502935, -2107570284, 638607502, 494230},{196608, 0, 128, 1140850688, -1255805332, 1228202, 1778384896, -2103957163, 486842, 1908032144, -1385400505, 1327811},{4288, 16777216, 0, 13641728, 935974144, -2099855849, 237139183, -667942906, -2096004058, -2096198223, 1303168849, 172071},{0, 17825792, 0, -1342177280, -600700158, -1164741470, 1897058917, 12, 1030144, -700730728, 464370309, 884439},{0, 0, 12288, 1075052544, -1220435380, 1031316, -1267204096, -2023227387, 995437570, 1616844176, 1434991453, 228959},{262144, 0, 8192, -2046820352, 1082266997, 2048350867, -835627339, -919766521, 1126235, 805306368, 1227905801, 1543709},{0, 68157440, 20864, 303431680, 397020781, -1252682217, -384413712, 1263836438, 1818068758, -417876247, -153260408, 10901},{0, 16777248, 0, 1174405120, 643113140, 1269205, 2091013488, 1073741831, 1510050, -1234157568, -2029490094, 1406291},{196608, 33554448, 16384, -2147483648, 1789785202, 1846713827, -964356004, 1481637914, 1742723, 1509949440, 113083671, 151322},{0, 48, 4096, 1881800704, -1811531763, 875180, -862616028, -1990172024, 1652779888, -211678936, 185430361, 732813},{327680, 68681744, 8192, 1901101056, 472789689, 611885, -1104041756, -1655582842, -725069238, 1001289077, -716927528, 321367},{0, 67108881, 134217728, 9470292, -381310208, 1029354, 1881447600, -1561329649, 577394, -1948778496, 1073741826, 1117643},{71680, 0, 16640, 17825792, 960055552, 2056674847, 1672097964, 128450584, 2052567125, -1425025104, 1794419332, 1691509},{6144, 67108864, 0, 805306368, 1364756841, 565349, -1747584112, 1542979592, 1806777, -1279747080, 1546387484, 994745},{262144, 48, 4096, -1073741824, 406241874, 2001894877, -826996308, 125335242, 207282869, -1595551531, -949940859, 533221},{196608, 83886080, 16640, 605290496, 1280881009, -1261409708, 1264849488, -884172605, 2056719478, -1825970532, -425952613, 1807031},{137216, 0, 0, -1709834240, 1790569290, -1990746973, 985200120, 1073741835, 1524168, 545381504, 144214344, 334466},{2048, 64, 12288, -1327454176, 398631429, 2035457495, 174699029, 20, 103936, 295960576, -719301998, 748397},{2048, 35127296, 0, -1610612736, -1255822307, 2073130542, -232086396, -2019178427, 2115667066, 1936996984, -1669332975, 503240},{262144, 48, 0, -1006632960, -1867999126, 796078, -70165232, 1073741841, -1759863855, 1850836244, -1989111215, 17489},{264384, 83886080, 8192, -1073741824, 607834237, 101929571, 1994895027, 292552722, 395596, -830877328, -2147483644, 953165},{0, 33554480, 4096, 805306368, -1213870846, 806466900, 237586800, 50075971, -204113289, 249024856, -1988848620, 1226517},{272512, 16777216, 0, 822116352, -599484343, -946946940, 773433298, -844103662, -624474807, 186122868, -744437818, 219977},{0, 16777216, 1744830464, 2654883, -1255805440, 1220076, -1111485836, 15, 1835008, -1356197220, -1073741797, 1126845},{0, 64, 0, -1036582912, -1464466819, 1006738, -327761568, 636485637, 1007843203, 1372904696, 29, 245760},{266240, 16777264, 0, 704643072, 1143249025, -649153723, -820845784, 397990235, -967665005, 1937474224, 1172320973, 1814107},{0, 17825792, 0, 1879048192, -431324411, 570330, 826889072, -1763081448, -644425473, -1218890008, 1419247619, 493261},{0, 16777216, 16652, 1896906752, -441101822, 1277420, -1546369260, 1244517463, 1960655984, 869522348, -155206967, 157233},{262208, 0, 0, 1900645952, -1673919988, 1421982, -357207706, 1530484103, 1489766632, 1237589053, 12, 1412096},{272384, 33554432, 4096, 719684128, 1208632217, 797947418, 989832744, 1096548381, 2139622451, 774834184, -1041484917, 1406562},{134217728, 16777280, 12288, 805306368, 649205897, -955737123, 2042436556, 945011989, 796442, 1665551800, -1805306408, 452438},{-2147483648, 0, 8192, 9459712, -130722048, 1151708, 271489788, 810905937, 404118, -1250949620, -2147483620, 1513007},{0, 16, 0, 1140850688, -1227958878, 966164, -327254016, -940572665, 1921807, -178793156, 1253922634, 584460},{0, 67108912, 20736, -1329528832, 1354011571, 1347603, -1849523268, 385613851, 1933883, 302028584, 2073147590, 398283},{0, 16, 0, -2046820352, -423288222, 1354902, -1442840576, 1197770119, -2049461491, 1619953892, -2007236601, 941198},{-2147221504, 16777249, 0, -268435456, -615432022, 955938, -1553331504, -1429209086, -627337281, 792777305, 28, 1511569},{65536, 50331648, 0, -1339523072, -425617380, -1307927598, 1400112468, 397769483, 1590131330, 1586075509, 1260690894, 1442167},{262144, 16777216, 0, 805306368, 1362477945, 705842577, 1656021672, 385700637, 1184032, -1418788864, -1762656249, 1546282},{0, 1048624, 4096, 722547744, -145829350, 1530514, -2065006592, 28, -354991616, -1971182388, 1518135132, 564168},{196608, 33554432, 0, -2113929216, 2067931204, 695123, 1112768512, 1161297946, -2059069307, 570722600, -2147483627, 1906771},{0, 67108864, 4480, 503316480, -517171031, 1329172, 1879048192, 11, -1925185536, -2095659100, 1882492103, 503422},{262144, 17825792, 12288, 587276288, -603596679, 991055174, 1406237344, 8, -648252357, 1917954373, -2146959351, 201689},{393216, 83886112, 16524, -1342177280, -331515743, 872450, -825749228, -1017311160, 1934935770, 256492248, 1960786635, 578173},{0, 33554496, 4096, 805306368, 75880625, -1693362721, 45501264, -1750313917, 801417752, 1517978376, 128743697, 620330},{0, 0, 8192, -1040187392, -330914966, 1277348, -239419392, -582132603, 897805, 1879048192, -1754154409, 1149904},{196608, 33554432, 4096, -737902592, 391837034, -2146263521, 39734393, 28, 177152, -570425344, 27, 1126912},{0, 1572928, 0, 1110048768, 910465170, 1400341, -451033032, -2009595887, 1842294638, -1032280344, -2147483645, 428163},{0, 50331713, 4096, 805306368, 1543690425, -67009019, -1747722968, -1423400755, -591027333, -1479257792, 231506583, 208659},{0, 67108912, 20484, 1881702400, 1196758137, 1199518, 1029032120, -1715732452, -2007927157, -1615488579, -1381856378, 433993},{-2013069312, 0, 0, -1320124416, -1213796755, 1220116, 1194922544, -348770531, 587681747, -1253404151, -731307180, 150854},{196608, 32, 0, 1879048192, -1152278267, 949410, -2032431892, -842998834, -833860075, -1909305920, -858246571, 1823963},{0, 16, 0, 67108864, -433411686, 1473242, 1027620864, -1073741804, 528195, -399538672, 1459728400, 211729},{131072, 16777216, 12288, -1837039616, 1764634026, -1395425763, -753938220, 1526756507, 899759, 1714559744, 52430100, 1408639},{0, 50331712, 0, -1340702720, -1071087013, 1158418, 685231224, -1684693888, -687469710, 666459024, -641627557, 243138},{0, 16777299, 16384, -972783616, -1227439475, 957588, 1555532656, -387414584, -649946409, 2128988004, 1281133845, 489177},{262144, 0, 268443648, -2046249902, -1180532405, 1963963732, 2003504124, 1073741826, 478324, 299273212, -1671380969, 1808342},{0, 524336, 0, 18927635, -1481260544, -174695086, 1774981412, -1858076643, -1643224106, 1586408228, 8, 205846},{6144, 32, 0, 1107296256, -442151579, 1548783084, -740640980, 1269599242, 1993608799, -1453865479, -1754441086, 1408095},{196608, 16777281, 0, -603979776, 1512126467, 1490083, 1135050752, 1688803287, -360107141, 2009635888, 1073741847, 730743},{266240, 83886128, 0, -254540416, -1213845835, -1391288812, 857825908, 1474320472, 2115476141, -277929191, -2095279786, 343173},{0, 67108896, 20480, 1892679680, 1279075225, 1413212, 335544320, 154140678, 947862, -1353938596, -1502058789, 461768},{4096, 16777264, 0, 8397920, -1195718144, 1023150, 982999040, -1654556603, 1594381972, 302045045, 3, 0},{327680, 16777216, 16652, 1879048192, 1161205849, 955478, 718985024, -578813946, 1615950537, -686729387, -1418318329, 405133},{6144, 33554432, 4096, 1879048192, 470177795, -1253147451, -1280628824, 355760003, -1870015121, 2003770124, -948406455, 1940400},{65536, 67108912, 0, -268009472, 289970186, -761889877, 1594776909, -1653483901, -195780789, -1223208616, -1664876516, 1358948},{0, 16777216, 0, 70975488, -147435076, 679122, -1372879088, -1073741801, 893022, 167772160, -2029518845, 371825},{0, 16777216, 0, -970293248, -1808142923, 546526370, -518126683, 6, 559027200, 1919517401, -960480617, 1815171},{65536, 0, 16768, 807927808, 1543911450, 1993757249, -1165393152, 23, 461863936, 780288768, 1747225027, 1104768},{0, 48, 0, 1150287872, -439270997, -829440980, 998808941, -1073741816, 450518, 0, 358910912, 1851830},{0, 84444736, 0, 1442840576, -81228375, 1097244, -1133656408, -1263983795, -727178573, -1696796349, 216559112, 1183964},{-2147418112, 1, 0, 1890615296, -1861396475, 1162640, -1143898112, -48758776, 1687384, 483249412, 5, 334848},{196608, 0, 256, 19922944, -1530330880, 420852456, -82259575, -963307262, 1876204765, 350013484, -191285359, 1193798},{67108864, 33554496, 20864, -1342177280, -599214837, 533254, -990658560, 1841460496, 226826972, 665845841, -414436861, 1907419},{-2147483648, 33, 0, -535429120, -71970478, 790009190, 1044054776, 2017722388, -1160308814, 2083036081, 410255373, 3515},{196608, 16777216, 8192, -1342177280, 1010128987, 1354689, -167772160, -2023176694, 1770167, 582013492, 1379139587, 1114923},{196608, 16, 0, 67502080, -144853334, 693778, 801591872, 201326620, 1690481, 1698042432, 342697044, 1492085},{0, 67633184, 0, -253427712, -804628468, 599586, -1275068416, 1239678981, 1540251314, -1562805048, 1170210834, 1124598},{0, 33554432, 16512, 1879361568, -716897515, 890663640, -119204767, -731906043, 2135292251, 1781678880, 542434653, 390848},{69632, 50331648, 0, -1342177280, 681648139, 1997513351, 1781693192, -1735131107, -1583674975, 652614125, 434999691, 590054},{262144, 17874944, 0, 1900101696, -172405492, 1486011818, -356845600, -1922251178, 822103100, 1851766622, -847249385, 247833},{-1945894912, 33554432, 0, 738197504, -1222185598, -460352428, 1050019404, 830629661, 1738691, -1353924008, 1313112078, 403485},{-2147483648, 0, 0, -335544320, -1732378107, 1219216, -708837376, 1976417627, 1565357, 1908260864, 23, 1836032},{0, 50331648, 0, 89128960, -1672560278, 679388, 271106048, 1137967122, 1028219399, 1858749288, -1844109242, 897078},{0, 35127312, 16384, 268435456, 1244960937, 823334, -778027008, -637009917, 2005497383, -1707202292, -2083152931, 1824384},{0, 1572928, 8192, 1107296256, -1255788989, 1027240, 1035550720, 1073741853, -696058937, 1446391809, 292141463, 1936341},{196608, 16777281, 0, 805797888, 352704585, -1122673495, 1723337664, 655656075, 521071, 244239308, 1073741851, 584892},{262144, 83886176, 4096, 1442840576, -516022103, 630996, 707641344, 23, 1807872, -1759625216, 48261659, 1359649},{67442688, 67, 8192, -301400064, 1549306228, 533354, 1602250620, -483491256, 2001267333, -1674657056, -2021886072, 1556014},{0, 33554432, 4096, -973078528, 1543854186, 19971, 2080374784, 432656149, 1185732, -338750148, -1073741818, 240539},{65536, 33554432, 402665472, 19989196, -427819008, 752274, 33554432, 1073741827, 1355229, 657956308, 498597896, 564843},{327808, 67633152, 0, -1324318720, -1853720413, -1757385180, -1411975794, 1229745986, 956636311, 2143564176, 59770837, 1907993},{0, 67108864, 128, 805306368, -1674014383, 1075328, 741065472, 29360131, 1879256112, -1961310536, 536870940, 451292},{137216, 0, 17028, 16785472, 927356672, -578135085, 450639656, -1921253347, 2039432569, 506593365, -1379464059, 343685},{-2147418112, 33, 0, -268435456, 1513472011, 1152417, -1827121080, -493354287, 909129, -1275068416, 3, 193536},{65536, 33554432, 0, -2046820352, 1756233835, 966235679, 376886668, 27, -930899941, 455826573, 359254235, 752985},{262144, 524288, 0, -1342177280, 836016133, 561305, 369098752, 17, 965837824, 2008757353, 24, 1119504},{69632, 0, 16768, 1879482400, -145143531, -946827818, 2061889488, 284950539, 376080, 820121796, 1846280209, 503514},{131072, 50331712, 0, 805306368, 1279301705, 948304, 332858228, 230963031, 764472251, 2008751468, 216911389, 1197788},{262144, 16, 12288, -267911168, 1630050413, 1209433, -1569226752, -660865011, 731026, 0, -1073741824, 1931145},{0, 33554432, 16524, 18251776, -1163570688, -690782820, 1646954708, -1073741804, 202950, 646774784, 2005055875, 540389},{196608, 17825792, 0, -1342177280, -1677019132, 1652657664, 176183161, -1803978853, 609884709, -286904763, 52962905, 1197107},{196608, 16, 16384, 805306368, 1264459865, -1018124134, -491568348, 1239991127, 2139343538, 605490772, -1907048253, 573373},{196608, 64, 8192, 821298720, 2067439761, -1672848793, -819919363, 387027668, 1607612123, 91313860, 432537618, 424544},{65536, 1, 12288, -1433370624, -147736948, -426549804, -676295060, -401820773, -2099804227, 138199520, 1137487130, 1836688},{0, 35127360, 4096, 823230464, -188101205, 1546924, -640252464, 2102460813, 1553012285, 1792749928, -2049703933, 1185740},{0, 0, 4096, 1141247552, -81146454, 1269294, 1501249536, 91750408, 584995, -784148556, -1073741813, 251825},{262144, 0, 12288, 1159725056, 818976938, 1473181, 2113929216, 201850893, 190660, 1394638848, 1122762781, 1809185},{65536, 67108864, 8192, 822083584, 1101412457, 955737, -2028448580, -725325813, 2005996831, 915333864, -1799271470, 771864},{268288, 16777296, 0, -1342177280, 17127564, -1668716541, 1394505497, 462946311, 787324, -1412458564, 3, 1808384},{0, 0, 0, 1507808, 357959936, 761005, -1409286144, -1942962348, 1294359, -1271116752, 6, 246784},{268288, 80, 0, 1898186464, -784821903, 1451520, -78089740, -1019917371, 391701, 1546900668, -904391157, 1929909},{0, 18350112, 0, 805306368, 382861323, -942760815, 807718352, -1946100468, -581052733, -472145148, 1284505606, 197853},{131072, 524288, 0, 1879048192, -1230681084, 963812, 1993933148, 1301282825, 1100022, -1827069952, 3, 205824},{262212, 50331648, 0, -1577058304, -1482510684, 418626962, 1647321903, -2147125623, -1411540520, -1766880524, -678864367, 194606},{0, 16, 0, -2046820352, 1543657541, 1083521, 0, -1073741824, 1547208, 2088189952, 28894741, 908925},{65536, 33554480, 0, 1073741824, 674884930, 609442467, -1097381535, -2089811965, 1104705350, -1961799423, -1016063535, 1286465},{0, 16777280, 8192, 1192263680, 1275156571, 157202, -1693464768, 120848387, 490259, -1912602624, -1864892388, 1413885},{0, 32, 0, 1478080, 2010568842, 679059, -600063952, 1190658050, 1149499, -1793523712, 17, 188416},{0, 35127296, 16384, 805306368, -1604806511, 1132650, -1938878128, 290485393, -1626237537, 249821349, -1073741810, 465820},{2048, 32, 0, 805306368, 1786943490, -158493917, 2010587928, 146901059, 365807245, 1973213629, -1073741812, 880917},{-2143223808, 100663362, 0, -2046820352, -1731022837, 1418894750, 448059308, 971957882, -976738696, -1631220320, 1265146440, 936153},{-2147483648, 65, 0, 67829760, 918962499, 637917, 0, -1492647936, -107199815, 286576992, -783477236, 1950171},{65536, 0, 384, 1140850688, -1255805373, -665403862, 2071008281, 337238103, 1497184, 19143928, 1913987206, 209738},{4288, 16777280, 20480, 1342177280, 646027337, 1967881109, 909273910, -1647201396, -679141858, 1471176145, 1550440398, 1908656},{0, 0, 128, -955207648, -615120302, 1532196324, -1262150507, 1465217933, 1143003, -1811939328, 814598556, 1690208},{65536, 1048624, 0, 1879048192, -1457066732, 1022684, 1845493760, -676046322, 593170240, 1044183837, -2147483637, 1323308},{0, 33554480, 0, -2113929216, -976833406, -2116830036, 339318873, -1738951854, -660770277, -558773859, -1653080051, 382643},{264192, 0, 20480, -1006632960, 807478131, -2049890779, -1229117723, 18, 1179648, -1987887104, 114918929, 753245},{196608, 16, 0, 1141506048, -456460628, 695258, 1107296256, 97255436, 240579, -1245822976, 1171807579, 1815998},{0, 0, 16520, 817954816, -1406887924, 1534700, -2057578792, -596115433, -673921065, -1183394071, 831221446, 377676},{0, 16777281, 384, 436207616, 1178900553, 768316048, 1635976028, 707626456, 1815420, 1914109952, 590886429, 1519484},{-2147483648, 17825793, 0, 805306368, 1706472475, 1021021, -241280764, 740556825, -917753234, -951358408, -638582781, 1695827},{-2147483648, 33554433, 0, -1342177280, 1512677652, 1489639, -104923136, 818732495, 1359417, 1580351488, 1097859083, 1832384},{0, 69747712, 0, -268435456, -1707457781, -996822384, -747137472, -2147483635, 812315844, 1176890838, 1550893458, 709081},{0, 0, 16512, -2044100608, 1143249002, -2100125654, -1672018299, -1737490409, -2028492519, -1857334887, 884030677, 1825502},{196608, 64, 0, -2147483648, -2128264787, -938385952, -79262256, 2, 897536, -579207168, -766747955, 620858},{-2147483648, 18350146, 8192, -637140992, 1758638162, -993018723, -1737271220, 947176528, -1093006719, -756600512, 283669575, 237328},{0, 16777280, 0, -1339817984, 1985291018, 876077, -1271954176, 540290691, 1921591, 506430048, 1104412692, 328783},{0, 64, 0, -2111467872, 1815773258, 1277413, 0, 443916416, 625536629, -576240868, 25, 202752},{0, 0, 8192, -950632448, -1806548716, 939564, 0, -1713373184, -1642480248, -1764288015, -662962159, 228039},{0, 67108881, 20864, 805306368, 956446731, 487095195, 1387676452, 1850267921, -1453722855, -287749024, -1557135358, 491427},{-2147352576, 66, 0, 0, 280306432, 1004705, -692085472, -332364088, 1809308, 1608239216, -1917549615, 552156},{0, 0, 0, -1040187392, 833995435, 2018949797, -383696708, -673447914, 48246, -598261760, 1086093399, 1553265},{0, 524288, 0, -2046820352, -2025151891, 678502, 1811939328, -969408506, 1708944486, 1662314100, 1073741841, 1863783},{2048, 0, 0, 70942720, 465655373, -494113641, -2025737871, -2147483619, 223714, -1731886232, -597164004, 1088519},{-2147483648, 33554449, 0, 805306368, -150595574, 1152274, -738197504, -199893667, 1954364, 130620856, 95158299, 1933257},{131072, 0, 4096, 1891663872, -1738996973, 1136092, -1212972608, -1073741811, 1529521, 2013265920, 1478769117, 1874586},{65536, 33554496, 12288, 805896192, -1404267407, 1971921730, -1222665452, -667346473, 433885003, 844978949, -2147483628, 1778281},{131072, 0, 17024, -2046820352, 1342789725, 1154566233, 1534301629, 1388386968, 1947972981, -732330652, 1951422853, 1121040},{0, 0, 128, 2523136, 2068226816, -2050011939, 1907640, -2096592445, 1537390, 364611752, -1145307114, 1598062},{131072, 18350080, 0, -1576648672, -421639507, 919830038, 842240388, -2090067748, 332499206, -1212259911, -1073741797, 1120531},{-2147483648, 1, 0, 68714496, -716000637, 1293228, -314321900, -1399324647, 1932910, -1787705860, 25, 1514820},{65536, 48, 16384, -2080374784, 400101547, 1220051, 1661048272, -2021654504, 1942710201, -797407355, 1005679568, 204342},{-2147418112, 33, 0, 0, -426878813, 1796584016, -223388555, 2005139481, 801501, 500776960, 12, 712704},{131072, 48, 0, 1107296256, 649240660, 766941, 121470976, -2147483620, 206446, -1336328192, -957846060, 1548392},{0, 83886144, 0, -973078528, -868826475, -1927987136, 1262585528, -595853300, 394199, 52711840, 148147270, 1935642},{-2147483648, 0, 0, 1879048192, 1369547274, 679001, 1150058496, -1462501364, 1602329, 9263656, 438931985, 783627},{0, 16777216, 256, 1174405120, 1732659371, 1530515, 1483980800, -2147483648, 1375887642, -566525347, -536870899, 1550150},{65536, 32, 0, 1882587136, 1498480658, 678811, 1982955520, -1073741800, 1131420, -1784738392, -1947205615, 1115354},{0, 50331712, 4096, 805306368, 1094828153, 1158683, 1893356684, 1302677709, 831658908, 2060274665, -2147483645, 329618},{0, 67108880, 8192, 805994496, 1278616338, -2096540776, -55256971, -1737490420, 1734194, -1965438556, -1031274479, 1145572},{0, 0, 0, 1140850688, -356179549, 1277348, 1833507420, -2062966072, 911860419, -106768051, 1516344644, 329033},{65536, 0, 12288, -1332707328, 1095057579, 2140323227, 1255098376, -2147483634, -540148608, -2072509064, 7, 748044},{0, 0, 384, 606635648, -189410493, 1465002, 1021762676, 6, 417792, 0, 536870912, 904156},{131072, 50331648, 0, -1332674560, 1479647491, 1162655, -1107296256, -1050818880, 1564426, 369098752, 23, 1144263},{262272, 16777216, 0, -2046820352, 1280612373, 1237419521, -563675693, 52256077, 1570173385, 1983058849, -707526650, 10569},{0, 50331664, 0, 1879048192, 738359298, 559235, 716331836, 1568244638, 223917, -895516672, 13, 1597440},{266240, 48, 4096, 823132160, -339145343, 1266642, -1814206652, -2147483627, 1948449, -1838563328, -1862008804, 1555057},{0, 67108912, 0, -1006632960, -800407228, 1123882, 0, 90778752, 241515, 2071281664, 9, 1230848},{65536, 68157520, 0, -1342177280, -598132726, 1166183936, 393697881, -166096101, -1144571111, 1196172037, -732089721, 152997},{262144, 524288, 8192, 805306368, 738883602, 886979, -83443308, -1073741822, -217988845, -1369853660, -2093149615, 1331992},{0, 0, 4096, 82870272, 886457202, 1935104685, 17729361, 17, 998768700, -1434397292, -684194360, 1818240},{0, 16777216, 0, -1339785216, 25604357, 752533, 1866893444, 1463584835, 986763384, 1057543277, 1073741841, 1431688},{131072, 16777216, 384, 436207616, -447294388, 1006702, -673841152, 13, 794624, 525472960, 721017239, 1328031},{0, 0, 12288, 605585408, -146693630, 1265066, 1275068416, 1518358993, 1762963880, 1061193448, 121110551, 1832725},{0, 0, 16524, 805634048, 1362401393, 1837205015, -713992431, 13, 1909234784, 680299997, -141856044, 1186500},{196608, 32, 0, -267976704, 952213787, 1331813, -1689583616, 1073741841, 1551250, 0, 0, 1321101},{0, 67633152, 256, 1882587136, 366087683, 1490271, 1641005960, 1132986370, -809256954, -1692784827, -1124072164, 579544},{137216, 67108880, 0, 0, 1275213824, 534058, 1326740680, 1507952652, 579353, 463643372, -1023909356, 783407},{0, 0, 12288, -1339424768, -180215549, 1203626, -1415816916, 17, 0, -1530033172, 1073741847, 1386199},{0, 67158016, 0, -1005027328, -461301612, 1465876, 747159552, 1123584579, -1974625072, -623201922, -2147483643, 747690},{2048, 80, 16384, 0, 1277534976, 446017688, -1898289915, -2025586668, 450606970, 1366951341, -2147483623, 383893},{0, 0, 16384, 1174405120, 282214978, 1027297, 1979711488, -938999784, 492751, -67108864, 133955596, 1502848},{0, 32, 128, 1882914816, -393635838, 1545178, 1677721600, 1379139590, 1121595301, 1435505729, 1715732506, 1729353},{0, 50331664, 0, -1339555840, -872007534, 390090242, 197608677, -814687416, -598868057, -408432292, 23, 807936},{196608, 0, 4352, 805306368, -662349819, -1211133032, -280439340, -949223395, -456755529, 1697761352, 922497666, 422631},{65536, 0, 8192, 1174405120, 733401365, -2045557795, 1789779321, 290222275, 654665, 2001277260, -1689963311, 1978034},{0, 0, 0, 1110770368, -340950357, 1021474, 341983232, 27, 1362944, -1602988852, -2147483631, 442484},{0, 0, 0, -2079682848, -1197080142, 957594, 1830027264, 1362362373, 1492297, -1795096576, 20, 1272832},{0, 64, 12288, 1140850688, -2133813173, 961560, 70156288, 1454374915, 886113144, -951725268, 20, 1779200},{-2147483648, 50331648, 8192, 805306368, -2004445180, 1207640, 1008537164, -1280514671, 1529433, 1464451072, 1419803348, 1340167},{0, 67108864, 128, 805306368, 1367461241, 1151145, -314191052, -1073741808, 92485, 507248640, -281483517, 1335205},{-2147483648, 524321, 0, 1879048192, 621360141, 1465563, -796453060, -1468792816, 1573994039, 640938141, 143130641, 1338684},{0, 50331648, 16512, 805306368, -1590296487, 1160552, -1781149332, -1073741795, 2081516804, 264865752, -1478897272, 937843},{262144, 83886128, 0, -325058560, -1865108965, 349466768, 982021297, 1194882060, 1523305, 1912602624, 8, 1316864},{196608, 32, 16384, 1107296256, -1138102621, 1084842, -1034794200, -1999265900, -1575672974, 1335855928, 387280588, 49805},{0, 16, 384, -268435456, 475944964, 1458311, 634753384, -1654279207, -698710250, 698522877, -44236268, 1135385},{0, 33554432, 0, -1072136192, 1506354002, 676756379, -1180744744, 1073741827, -993243966, -569991936, 64225293, 1701970},{65536, 65, 0, 805699584, -1152005523, 1023138, -1227210752, -1505230828, 1293718434, -332429787, -724566005, 1700251},{0, 0, 4480, 1155563520, -1807863645, 703914, -1952955448, -1065615357, 842811, 1958234208, -104286131, 1901338},{0, 0, 0, 1175879680, -1056843710, 693226, -1648508928, 13, 875520, -667828224, 1073741851, 1363593},{0, 16777216, 0, 67108864, 724213860, 750435, -1275068416, 5, 1651712, -1424408576, -1073741801, 1549733},{196608, 67108864, 8192, 1879048192, -1674537709, 2144632896, 1786791944, 11, 1950918144, -1098855163, 1444675611, 209780},{0, 1048640, 0, 805306368, 28612609, 565331, 1610612736, 1416364052, 1149840, -1348245540, 125646225, 411773},{65536, 0, 0, -973078528, 1342554805, 611291, -19185664, -1073741811, 1772715, 1621953228, -2147483631, 1024197},{196608, 67141648, 0, 1879048192, -1492576244, 1334418, 1987543040, -881032058, 916084356, -1958467981, -942669817, 1348733},{0, 68681760, 0, 1073741824, 1278280106, 953184, 872415232, 11, 1736644, -68965740, 1413480458, 1932619},{65536, 33554496, 0, -268435456, -242861932, 698960, 2131842608, -291151029, 1669786340, 846499493, 3, 404598},{-2147221504, 0, 0, 805306368, 295999569, 30699665, 720585960, 981205396, 1134409, 631768272, 77332497, 7245},{65536, 0, 8192, 1882619904, -1727981547, 1291228, -1562620808, -1917215215, 1363503, -2135635580, -1712016168, 1776176},{-2147346432, 64, 0, 1073741824, 1003146597, 611217, -1686789164, 1955652805, 157513, 472514560, 64487427, 1265785},{262144, 35127296, 0, 1107296256, -984951476, 750438, -1753714384, 1340618769, 26276086, 1580540800, -785121260, 1335603},{131072, 48, 0, 805306368, -2134040549, 1461086884, 1046087064, -2147483631, 212664, -1313993848, 1222639632, 1102983},{-2147483648, 33, 0, 1342177280, 625090818, 949485, 1580799872, 1033226516, 246503, -2080374784, 1468360513, 1907769},{196608, 16777280, 0, 807698432, 2057404521, 939117, 1058672956, -2031545129, 330562, 1845493760, -1858009196, 1356913},{262144, 33554432, 4096, 805306368, -993369334, 630610602, -2028541740, 7, 897800192, -613329156, -886267257, 1925714},{0, 0, 12288, 1140850688, 274088346, 1464977, -642514944, 21, 1432576, 671088640, -2147483625, 1146745},{0, 16, 0, -1070923776, -511362990, 1031194, 1958972168, 24, 1702400, 1811939328, 0, 244736},{264384, 83886080, 8192, 1879048192, 1280356357, -1626593774, -15287757, -949109290, 857564797, -616115107, 467140629, 1924734},{0, 65, 20608, 805306368, 1544206513, 549096, -637534208, -107709373, 2106254020, -925449280, -1384376615, 1599391},{0, 16, 8192, 3899392, 616164608, 1267235, -733233152, -2066481148, 895933, -762740736, 225295444, 1365722},{0, 0, 0, -1040187392, 556376946, 1023513, -671088640, 1301595715, -632187843, -2022029864, -2147483637, 1681449},{71680, 0, 0, -1006632960, -1610237814, 1223954, -1506592892, 1526489160, -1345843947, 555044553, 1073741846, 1542508},{0, 16777216, 12288, 807927808, -1707753462, 1219554, 1952876720, 6, 569344, 1719473088, 342622234, 1159801},{0, 0, 8192, 806882816, 959828227, 1460767, -1409286144, 1254928592, 901328, 1185988608, 1073741847, 920343},{0, 0, 16768, 738197504, -1867923327, 1353882, 1350929284, 8, 1350840, -2071576576, 1941962763, 560038},{65536, 0, 0, -267845632, 293976076, 1506386081, 259397481, -2147483621, 393590, -1723596800, -1073741801, 1934798},{0, 0, 256, 1174405120, -1601529715, 1137470880, 1298353829, 6, 1098907648, -789952671, 536870932, 515768},{0, 32, 16384, 808878080, -1867474772, 1162640, 872415232, -1877475311, 1357392, 474619412, -1610612736, 1519283},{-2147483648, 17, 16384, 688128, 1096677376, 882073, -1600615656, -1379618419, 960433, 160530432, -914620413, 1322910},{0, 67141632, 0, 806748160, 562149489, 167465, -844857344, -844103673, -573270648, 38615682, 441245213, 1274085},{0, 0, 16384, 1882587136, 1092985093, 1267109, -466092032, -1073741809, 1043457, 1329992512, 1073741835, 196367},{0, 0, 384, 67108864, 356581709, 1020651, -1263337472, 174325780, 1098931, -732296988, 884294352, 252468},{0, 0, 4480, 1778384896, -427419644, 630918, 2016559104, 25703191, 230244, 0, 1029447005, 1128262},{0, 0, 12288, -1340702720, -1171127805, 1152340, -2080123796, 1417689155, 756555, -1590916252, 1247626516, 1762998},{0, 32, 128, -1342177280, -1043187700, 1400020, 765607936, 1512411274, 1940337, 615694948, 2046296069, 1541689},{0, 16777216, 268, 1494253568, -1488014189, 748946, 2098630692, 377845719, 395782517, -1217063347, 1901551060, 1131290},{0, 0, 0, -1340571648, -1053392125, 72523092, 1891943304, 4718592, 71522873, -1128920520, -882899645, 1603760},{196608, 0, 4096, 526688, 684577792, 1863693275, 1719519108, 29, 1158144, 1303379968, -1851523065, 1547889},{0, 0, 1207959552, 1313443, -1196831387, 1539244, -1199800320, 25, 1689624, 2084329408, 13, 1552469},{262144, 33554432, 0, 805306368, 1622227049, 1502264363, 1269126997, 7, -1261860864, 1871776616, 1515811732, 1827404},{0, 0, 0, 1176895488, 1082308716, 543649, -1780465664, 1518985293, 514938, -2013265920, -998652390, 390343},{6144, 16777216, 8192, 1879048192, 123054594, 769439, -675416120, -612270972, 719019, -1565566076, 461658125, 568045},{65536, 0, 12288, 1073741824, -1455095134, -2024579752, -629337144, -1073741821, 498826, 1820819456, -2147483628, 1731175},{0, 17, 384, 1879048192, 657862674, 1269141, -1064662184, 1834792333, 1769237, 1955187216, -1329296751, 1543029},{196608, 64, 0, 805601280, 1633455497, 1409113, -1296558116, -933232632, 554629, 0, 1474320320, 547000},{0, 50331648, 8192, -2113929216, -625917788, 1275286, -256189476, -2147483620, 1546425, 332944804, 27, 1774526},{2048, 33554432, 0, -1342177280, -1940511924, 1464964, -2025201664, 1526489227, 959922, -2106173576, -679910837, 1327426},{6144, 64, 0, -1332016640, 1280612355, 893026, 1803091232, 1256194071, 580170, 414679040, -1073741794, 1130760},{65536, 0, 0, 1140850688, 952213570, 678821, -745350396, 1073741844, 623024, -307200000, -2009071591, 539056},{0, 32, 0, -2046820352, -1869989787, 890384, -378103840, -1073741817, 316233, -2026107312, 1474582810, 1542490},{2240, 67108864, 0, 805306368, -1498242556, 256984466, 450653039, 17039371, 268625935, -164232956, 17042457, 1045558},{0, 0, 128, 100663296, -1807375755, 806771370, 1772225288, -1709076918, 1102990, -1275068416, -348906156, 910244},{196608, 16777216, 8192, 0, 388369850, 1006741, -2113929216, 3, 156672, 1674972756, -1752864876, 1132082},{6144, 0, 16384, 338167168, 982398981, 1175936421, 850965233, 11, 1218087936, -1992975732, -2143027180, 1153592},{196608, 67108864, 20480, 1880522752, 2712177, -523360749, -1431204371, -569638909, -958853922, 329288064, -1073741816, 529356},{131072, 16777216, 0, -1845493760, 1641914386, 382630937, -2022369655, -2147483645, 408174915, 1728398188, 11, 224571},{6144, 67108864, 0, -2078900224, -83748693, -703443486, 641088081, 493932954, 245133, -740864512, -1705713654, 31748},{131072, 16, 0, 1073741824, -150547013, 1133584, 2137243648, -882638825, 1528436, 1152794624, 7, 1481894},{262144, 33554448, 0, 100958208, 1994009218, 760741, 1134335924, 1129316756, 234044, 1650114592, 1073741835, 102402},{196608, 67108864, 4096, 805306368, 1279623745, 871594, 57955896, 27, -1584288256, 978098452, -1073741802, 516789},{266240, 0, 0, -266698752, -801601132, -871284500, 511556725, 0, -574619648, -1731378051, 13, 1956864},{0, 64, 8576, -2147483648, -333061715, 1384345092, 1300944173, 1535451994, 199343, -776856804, -1169075510, 1727053},{0, 17, 0, -1342177280, -779757563, 572376, 101712800, -1482420194, 1739642, 1630814896, -2133837228, 513159},{6144, 16777216, 0, 86016000, 2069015179, 1989057367, -887787308, 240910359, 1144038, -2037741036, -1073741797, 902358},{262144, 0, 12288, 1109688320, -1432207261, 1471206, -1561985024, 5, 502784, -1000865792, 1315176468, 571218},{0, 0, 0, -1340702720, 1629561603, 1227873, 1518190592, -2147483637, 1934799, -461864960, 7, 752640},{-2013265920, 64, 384, 805306368, 1275181129, 1409688, -585449472, 730232469, 412399289, -515632723, -1238832491, 1565368},{201588736, 17, 0, 805306368, 268769298, 1403681, 396172044, 2005850775, 761531, 1073741824, 17, 1088512},{-2147352576, 67108944, 0, 1479966720, -1408603231, 949568, -1483188248, 2045555598, 1433522, 796371664, -975175657, 540030},{397312, 67108912, 20480, -1342177280, 1546715569, 1016407590, 239940765, 133203915, -518118683, 2058872961, 504483288, 807560},{0, 16777216, 0, -2046820352, 1359026331, 1462885, 117407744, 27, -2118061056, 192517932, -832045029, 1112441},{0, 0, 16388, -2046820352, 928703116, 678867, -793722880, -1955069948, 197706, 875367292, 2005575435, 885630},{0, 17825792, 0, 805306368, -459103476, 687642, 2104688640, -1758461929, 1694565938, 104211081, -1073741823, 937056},{65536, 0, 8576, 1073741824, 470641795, -577590359, 591058024, 26, 0, -1674018744, 1843451924, 757427},{0, 0, 12288, -1006632960, -1941585501, 1199424, 885456896, 432799755, 693709, 1509949440, 14, 940544},{0, 67108864, 12288, -1711276032, 1356505627, 1530521, 969834496, 194023124, -568684740, 2065125573, -572522490, 232120},{2176, 0, 0, -1342177280, 1543649300, -686522173, 249494071, 464781342, -636644929, -1447109784, 1542717463, 1830106},{131072, 16777216, 0, -2046820352, 961683563, 1292544979, 1383384905, -2147483625, 1738183761, 1857423932, 1073741827, 1458509},{333824, 0, 16640, 1880850432, 77712737, 1511101087, -1707351100, 1075840983, 968988027, 48696928, 1736194318, 1827749},{196608, 0, 0, -2079064064, -189415251, -1575973330, -1633495487, -2147483626, 1691022, 1543503872, 1073741835, 1526179},{0, 48, 0, -1037500416, -1495662451, 760796, -1140850688, 62920131, 218696, 1842118656, 13, 892928},{65536, 0, 0, 805306368, 1361232652, -774403495, 1722766400, 26, -535243552, -626125524, 1073741828, 1729957},{131072, 0, 12288, 1879048192, -1064683517, 1350800, -1979711488, 26, 977449984, -562211644, -719060963, 1974906},{0, 0, 8192, -1340669952, 72721157, 1031251, 1543503872, 14, 486871, 601522176, -2147483621, 1725401},{329728, 67108912, 0, 1879048192, 1543638865, 1758283932, -1240451247, 1579998356, -950767796, -605893192, 1556873232, 239477},{65536, 33554480, 16384, 805306368, 1278515337, 1343506, 2010662768, 245891089, 748501, -945336664, 126877709, 1926782},{131072, 48, 0, 1605632, -1453659904, -762413862, -417768472, -605440489, 1386266, 890980020, 238361422, 943966},{266432, 0, 0, -2147483648, 280270922, -1651592021, 179956663, -718690918, 928071946, -1317840296, -2089539891, 1521041},{0, 16777216, 8192, 1077182464, 992668813, 750437, -329365584, 1073741849, 1676518, -1951361044, 1315176471, 961156},{-2147483648, 65, 0, 1141605760, -1717416572, 678876, -2145910784, 1745913876, 19377, 1413333956, 1389101070, 1892680},{196608, 0, 0, 1543503872, 11870725, 701545, 1041239724, -2011108661, 1048953, -126271488, 1073741840, 1568269},{0, 67125248, 8192, 825262080, -1531821310, -1349604504, 2016434833, -1015539573, 920292424, -807327614, -620997735, 1352238},{0, 0, 0, -1340571648, 22356740, 1273241, 741310464, 3, 1855566, 1784743116, 14, 320512},{65536, 33554432, 0, 1175060480, 960640682, 1530527, -637534208, -731009148, 1300701, 934248448, 1160773643, 1351865},{2048, 50331712, 0, 805306368, 1359067265, -858688983, 853912228, -1859585961, -1554282785, -2032168663, -1717043177, 735651},{0, 68681728, 0, 805863424, 13238857, 873681, 0, 0, 1144271, 2050538736, -791150584, 1326396},{266240, 0, 4480, -2147483648, 959902021, 1301238365, -1411253268, 1302443720, -1185437256, -666051539, -536870908, 914339},{0, 16, 0, 1879048192, -1585326076, 542880, 0, -885784576, 758353, -474870988, 1249116189, 479562},{0, 33554432, 0, -264763840, -606461932, 949784, -1134864736, 3, 0, -298248316, -1752694757, 90491},{0, 32, 16512, 808714240, 473208905, 1154372737, -1766435152, 1371042522, 747177, 1427914752, 1682967511, 1328973},{0, 16777216, 0, 0, -2128174230, 185512616, -1866970968, 492830733, 758231, 1926890572, 1073741838, 282071},{0, 0, 384, -2080374784, -1252646555, 1775410030, -1338392108, 24, 608410907, -1320299303, -352738031, 1718182},{-2147483648, 1, 8192, 33554432, 2002178157, 395416145, -662912328, -188466617, 246750, 901480448, -2123250852, 1740311},{196608, 0, 0, 35979264, 2026034525, -825328807, 601296428, -2038373669, 918489, 1882620028, 1423789379, 942199},{0, 33554432, 12288, -1508311040, -1412259819, 748306, 1879048192, 296486851, 899533, -1506377728, -776922749, 1387207},{0, 33554432, 0, 1075351200, 2066631234, -535989465, -528693384, 506462215, 1733856, -1344077824, 1557921821, 1935570},{0, 16, 8192, 1879048192, -1254023156, -489841372, 1614004277, -2147483621, 1978302, -1177731072, 1580204038, 1529395},{0, 0, 0, -1340864000, -1680694523, 873634, 1214332928, -651410300, 961362, 402653184, -1073741818, 41057},{71680, 1048576, 0, 805306368, 1786878093, 1415015059, -350553672, -985546213, 1567838, -1226605536, 1532755985, 1699924},{196608, 67141648, 0, -1342177280, -1979041780, 416066150, 1109298728, 1210376849, 1020943077, 1983346486, -1049624547, 841752},{131072, 68681728, 0, 1610612736, 732086556, 1896764627, 318868781, -2130386021, -481401073, 1132390300, -1763966954, 962929},{0, 48, 16512, 1073741824, -1958329731, 611814, -102739796, 1363148802, 1974215, 487866368, 1661490142, 10056},{0, 48, 0, -1876361216, 1774625027, 1528415, -1370612708, 1474058126, 945022, 1409286144, -712392165, 208945},{131072, 16, 0, -268435456, 371884802, 34780011, -1838103680, 26, 227840, 1360314368, -2088501231, 1769280},{262144, 50331680, 0, 805994496, 950083921, -1554619675, 789745545, -2010906603, 1530598, 1525088256, 1073741852, 1690829},{131072, 18350080, 0, 1879048192, 1443182610, -959006053, 1866305909, 20, -811926563, -1564888003, -1073741804, 1108446},{0, 50331665, 0, 1879048192, 1792868370, 1151811, -373931684, -1529235045, 1125087, 974526628, -1073741813, 1730980},{262144, 32, 0, -973078528, 1348010259, 1901181533, -968336331, 1529085972, 1958851, 495681536, 438042650, 1740220},{0, 0, 8192, -266797056, 1817355012, 619035, 0, 397934592, 1846844, 1893580800, -2048393215, 1832864},{0, 67108865, 12288, 1107296256, 2084910661, 1967811365, -2056646372, -1419402038, 735154, -475742208, 1361152661, 1354613},{327680, 50331712, 0, 1879048192, 1279869545, 890331218, -1277748420, 494155021, 26861274, -1632035484, -1950613501, 1542667},{0, 0, 4096, 1174405120, 1967817293, 875757, -660062208, 1, -1282722816, -948268624, 17, 283242},{0, 16777280, -1476395008, 807833120, 1761949777, 1277405, 1275068416, -877362040, 557753, 1310170044, -1073741820, 515204},{131072, 16, 16768, 1879048192, 1275762802, 1092570, -1642741760, -2090336253, 1158787703, -555348732, 1682967572, 1548198},{0, 67108912, 0, 807667104, -331048815, 630016, -1387867132, -1016579823, 386115277, 2143511452, 342884363, 900118},{65536, 0, 8192, 1073741824, 293984405, 678875, 774160384, -2086666226, 1724812, 1345978368, -2014982630, 1367762},{0, 0, 16768, 1075445760, -148757870, 1421990, -399785984, 1135098459, 19894, 902660096, -1610612733, 910307},{-2147418112, 1, 0, -266010624, 402995202, -1311920999, 56169668, 639179534, 1979115, -984757832, -887095279, 435533},{0, 0, 256, 0, 13771520, 1289369, -387530752, 16, 946176, -241384124, -1151279591, 1979163},{264384, 32, 20480, 1879638016, 1724714005, -443059565, -1438336414, -1684235113, -1252575618, -1930732640, 1537258817, 894699},{-2147483648, 67108865, 0, 806813696, -788440927, -959095784, -125116887, -391257264, -2024004738, 1393088236, 7, 1512448},{65536, 50331680, 0, 24183168, 656813312, 759929813, 736153921, -1806696434, 1158568879, -567239471, 1073741827, 341260},{0, 16, 12288, -2147483648, -86924733, 1490148, 968132176, 344009884, 1313749834, 827923497, 92360259, 963454},{0, 0, 0, 1076264960, -2116697678, 1031330, 337936384, -1073741817, 1133628, -603979776, -2147483645, 1367042},{0, 64, 0, -2111435360, 1514828106, 766941, -1334509568, 1526726668, 719583, -320906472, -812646371, 1843986},{131072, 50331648, 16384, 1879048192, 1084266498, 1157921, -1545797632, 477419796, -598459120, 1933610440, 1903689748, 1362488},{329728, 1572864, 16640, 1879048192, 1216694625, -1504531557, 1997716529, 1073741853, -1472110149, 1927331225, -1141531442, 1941411},{196608, 0, 0, -2147483648, -794156372, 1022880, -344817664, -1073741795, 1711499, 738197504, 23, 1518592},{327680, 67108864, 0, -1071315456, 1549411258, -1592908258, 2004583917, -889609958, 908720, -1978017272, 87556125, 248241},{69632, 0, 12288, 805306368, 1543837707, 1971358723, 667118244, 1511522331, 1529251, 529121280, -1765539814, 1744566},{0, 0, 0, -2078863872, 614572205, 1267171, 1232535552, -680525820, 1926145, -469762048, 1073741845, 42420},{0, 0, 4096, -268435456, 1631666957, 1207379, -253997648, -1796970476, 1724282, 1367098712, 162102347, 1122997},{0, 50331648, 0, 1879048192, -2126438140, -1395497624, 1405307752, -2147483645, 1612054710, -1031483859, -857120693, 1819874},{268288, 0, 8192, -1743224832, -422939574, -1189759466, 119219048, -973033151, 1556859, 984697096, 195069323, 238103},{0, 33554480, 0, 33980416, -173715798, 1162656, -1741255880, 3, 386644480, -1575252628, -1968701429, 902323},{0, 16, 16640, 1174405120, 677210802, 881891, 2024751104, -1857245679, 1905156984, 1405982572, -1104061436, 321251},{0, 0, 0, -973078528, -794705237, 611752, 881530684, 3, -1538752162, 1821054809, 1073741825, 1339987},{-2013265920, 0, 0, 1174405120, -96898733, 1416740, -249706876, 772447174, 238501, 536870912, 299892747, 1161644},{0, 1, 0, 33554432, 389888163, 886125, 671088640, -101652978, -842814530, 1491537464, 126877723, 1695170},{268288, 16777216, 0, 805306368, 1090677833, 1421969, -613031864, 1078568516, 81502408, -562098652, 1515031124, 729826},{0, 0, 12288, 67108864, -1496776373, 1342374, 0, -596342912, 947055, -1653522432, -567541744, 1109775},{0, 557056, 0, 1895858176, 665202195, 679149, -716895308, 16, -1623195648, 1471819447, -1073741813, 1131821},{65536, 0, 0, -268435456, 296370188, 614555, -1347877672, -1073741816, 1565025, -782123008, 1520263698, 363848},{65536, 84934720, 24576, 805306368, -1702496079, 365469888, 708626236, 638858075, 1359713093, -1478363939, -783199987, 1930789},{65536, 0, 0, 67108864, 1698759499, 2089904875, 987709485, -1073741796, 1119293, -432324608, -1748215084, 1775819},{327680, 68681728, 0, -2111373312, 668278869, 1293847, 2068037632, 1174667265, 1984808310, -566559267, -1918631929, 1317324},{0, 50331664, 8192, 1778384896, 1755447306, 337074843, 1165791557, -1702517557, 206436313, -209877587, -884436963, 1126282},{0, 33554432, 16384, -2147483648, -2135350398, 1758434410, 495715456, -963641318, 221255, 2053685248, -2108405743, 1159733},{0, 68157440, 0, 1174963776, -422483302, 1539498, 0, 102498304, 247836, -406608352, 1161560071, 1555551},{196608, 33554432, 4096, 1744830464, -651866107, 757166, 799113216, -1073741797, 626663239, 710186109, 1162678363, 1780618},{0, 0, 16512, 469762048, -1853794159, 34637968, 303062372, -2147483622, 1851822, 1370390528, 537395204, 401329},{266240, 16777264, 0, -268435456, -1875604966, 38698090, 1198876244, 435264965, -405715326, 1800290340, 1316749323, 903170},{272384, 0, 12288, -268435456, 1356464669, 1611486297, 1511585651, -2021654514, 642468, 1436850308, -829888693, 218830},{0, 18350080, 0, -2080112640, 398014317, 1220117, 335544320, 1073741850, -1865706472, -961206116, -1736703977, 224673},{262144, 33554432, 12288, 1880850432, -390987758, 758426, 181993472, -1073741821, 114742, 786189112, -1047483442, 1849913},{-2145386496, 66, 0, 1174405120, -519964604, -682339744, 1897187129, 722959415, 209753, -387953348, 1073741845, 719072},{0, 0, 0, -1073741824, 1363493746, 622683, 942867244, 1073741827, 113013, -977043456, 50069526, 1849790},{196608, 0, 0, -268173312, -1051279075, 365523816, 916193636, 30, 729088, -536870912, -2147483631, 429337},{0, 33554432, 0, 33554432, -1764621429, 18240848, -1281418204, -1650720760, -905026086, 1786626065, -1023138534, 4144},{0, 69747712, 384, 1879048192, -2040858614, 175104, 1838172256, 1214251022, -1304800122, -166301242, -531857125, 1172396},{0, 0, 0, 1110085312, -1262938237, 1211476, -1065663928, 1316487173, -409529252, 990892208, -1012924402, 377914},{0, 84934704, 16384, -267059200, 1547870234, 1479784, -2048844576, 1578106887, -414271769, -488475936, -812300979, 1707794},{0, 50331680, 0, -2145910784, 1220457067, -414535087, -513686504, 1142685719, 2052994888, -1235680228, -2147483640, 1240295},{65536, 33554432, 12288, -1778384896, 1218789387, 1226079, 1382121472, -2147483628, -497741624, 780471864, 40142171, 768573},{0, 0, 16512, 101351424, 1766957706, 1538653, -67108864, -616824803, 351711, -1115923852, -302407476, 1552297},{262144, 18350080, 0, 369098752, -1593397143, 1018770, 1323188224, -2046172344, -859620542, 320159277, -1914141675, 1327324},{196608, 33554448, 0, 0, -1139963284, 1152284, -161562624, 416022541, 253861, 461160448, 1356333083, 591124},{0, 0, 8192, -1338736640, -106815228, 1399452, 484526124, -930815666, -2007537951, 1481115784, -963590717, 1961509},{0, 0, 8192, -2147483648, -1942576822, 1151172, 497211380, 1573388294, 1664084, -910999552, -634290275, 740218},{196608, 0, 0, 1142227360, -146443166, 1291620, 503316480, -670826470, -2142943209, -114982527, 95420440, 1713175},{0, 17825792, 0, 1882849280, 366348810, 344747181, -875111184, 3, 83968, -1012686520, 23, 0},{196608, 0, 0, 1881669632, -1759411965, -1559276382, 1260575217, 1512674001, 1342978, 404835812, -1914404222, 1371169},{67108864, 50331712, 0, 805306368, -335087604, 1421442, 495730688, -1538129894, 2023465902, 1454706292, 1513619459, 634074},{0, 16777216, 0, 1177060032, -701927867, 1220050, -1720024044, 68419595, 2080959868, 2117517705, 14, 267264},{0, 16, 12288, 1879048192, -2126913510, 1354394, 1823261536, 1100264323, 1723100, -1540014080, -2147483635, 933378},{0, 0, 256, -2046820352, 1490157931, 1197471, -2080374784, 451411991, 918740, -999023892, -246415146, 1710771},{0, 64, 0, 1174405120, -1059962211, 871842, -1049280512, -1704984575, -1508581523, -1614855375, -1073741821, 212373},{196608, 0, 0, 1610612736, -1062624764, 1203112, 1004182132, 30, 1171456, 102123152, 1073741838, 92590},{0, 16777216, 0, 1174863872, 1090893996, -485536623, -1662825168, 1311768605, -884993821, 976241237, 28, 856064},{272384, 16777216, 12288, -1342177280, -397109171, 545810562, -1683458955, -929266211, -1819597915, -476489123, 1214597009, 1166246},{0, 50331648, 0, -1071120384, -1951022685, -271469212, -788295232, 1371537409, 328269068, 1918649245, 14, 1128448},{65536, 0, 12288, 1141178368, 1975120203, 1220141, 1927807864, 1173618702, 1930330151, -121650315, 28, 965491},{0, 32, 0, 1474560, 1472340853, -443368047, 95487004, 20, 948967, -1595473920, 1142947860, 1565785},{0, 33554448, 12288, 805306368, 457291011, 1359582173, 305955281, 379846686, 947845, 1205813248, 502530065, 1332834},{262144, 16, 0, 815847456, -1858960471, 2072886352, -877392264, 1316534861, 270247, 280641536, 192710427, 949169},{0, 32, 16384, 809009152, 1619605393, 684907, -2013265920, -729206956, 777327586, 994319569, 1416709454, 1443460},{0, 0, 8576, 1880653824, -1177881083, 611098, -33554432, -1073741795, 1559965, 0, -348364992, 916348},{196608, 0, 0, 1881571328, -179977982, -1470980842, -1970781219, 23, 219136, -1072244068, 1211476419, 911910},{268288, 0, 128, 805306368, 470063185, 1418745985, -82544280, 10, -870631424, 830443016, -302514150, 1731254},{4096, 0, 0, -1340440576, -616488190, 395033496, 383902076, -2147483634, 1637795, 629669888, -2147483622, 374177},{196608, 0, 4352, 805306368, 1711729924, 686981, -1038761984, -2124677097, 1952719, 0, 1030755840, 1571747},{196608, 0, 17024, 805306368, 22733058, 617561, 2135703552, -1914380780, 1574433, 738197504, -1261928504, 1701826},{65536, 67108864, 0, 1174405120, 738550285, 690179, 1390526464, 433848324, 947398, 1320583168, 0, 703609},{6144, 17825792, 16384, -451903488, 1544378522, 2080531975, 860826525, -1706456934, 1326158246, 450782233, -1796134782, 1514049},{0, 0, 0, -1342177280, -1856625916, 868448, -996386008, 29405709, 897079, 0, 1073741824, 1719199},{0, 50331664, 16384, 24164361, 953811456, 678885, 383798596, -2025581116, 1557357, 1930756096, -2147483645, 1450872},{0, 0, 0, 1174405120, 12993181, 1461801, 1668193040, 3, 0, 1006632960, -1755840509, 120258},{0, 48, 0, -268435456, 554620164, -838236069, -1601888719, 1268776971, -1966209431, -300513184, 1073741850, 568803},{0, 67108865, 0, 805306368, -1674927183, 802884, 73990144, -1534853117, 1767531459, -902898488, 1073741837, 1941576},{-2147483648, 17, 8192, 1879474176, 1472844812, 1489489, -1525399552, 1713399705, 1172398, 1695825920, 1357381658, 1945186},{327744, 64, 0, 503316480, -509300055, 265578640, -2099024333, 288931012, 430650, -658716600, 16, 152836},{0, 67108896, 128, 805306368, 1103661465, 873817, -396387744, 489947138, 1728422, 601505792, -1552312826, 567111},{0, 16777216, 16384, 1677721600, -1052441846, -485657362, -1025041624, 17, 1262854144, 998136484, -1927959983, 347875},{131072, 0, 12288, 1879048192, -1154842363, 890402, -2092610824, 1527513102, 1649694129, 842859116, 23, 1974064},{134486016, 80, 0, 1901068288, -1531575887, -527729746, 665955236, 883079424, 1436153575, 1960761340, -1073741816, 809343},{131072, 48, 0, -268435456, -1699364589, -401427360, 316444292, 26214421, 1485504, -146701932, 29, 94208},{131072, 1572880, 0, 738197504, -1954383861, -636912742, 2052808229, 1570766862, -1286887521, 333478505, -1660682213, 1560034},{-2147483648, 33, 4096, 1879048192, 453949451, -267238481, -1977871936, -495698796, 1980128, -536870912, -775684083, 1339957},{0, 35127296, 0, 1107296256, -190668684, 1201644, -469762048, -1839612325, 718942433, 1924410905, -1680605173, 1667203},{268288, 0, 0, 805306368, 558801179, 1489555, 853795092, 3, 176231424, -1617340128, 438853018, 1717272},{0, 557056, 12288, 536870912, 741945610, 1266975, -1519085992, -2147483622, -685944751, 195246075, 447313102, 1954327},{262144, 0, 12288, -266043392, -794181606, 1080720, 308019200, 1073741824, 1367474, -796753920, 1529442693, 1575646},{0, 65, 4096, 1174405120, 356384778, 1422057, 1021165568, 2046091022, 550469, 954138624, -2018719462, 284391},{0, 64, 4096, 1174405120, 20101195, 1137283, 261279288, -1910767602, 378789, -1580970916, -1004797941, 1373992},{0, 0, 0, -2046820352, -1596808604, 875730, 1787124232, -920649717, 952551, 1409286144, -1073741816, 903306},{327680, 0, 16640, -1329528832, 1350645866, 1209763, 527335424, 4, -1362014208, -207071351, 659297812, 271034},{137216, 0, 16384, 806617088, 1250089033, -527330280, 1924381753, -2147483645, 212448, 566837248, -484645669, 546738},{131072, 48, 16384, -268435456, 1346453882, -1542642147, 106695468, -886308850, 1765234, 1708103496, 8, 1735168},{0, 33554496, 12288, -266665984, -1607428070, 1142240, -988050440, 245659217, -355187763, 1541014660, -2097387177, 1775152},{131072, 18350080, 0, 1879048192, 1460246531, -728580701, -1570632188, 502126091, 823215376, -1356925811, -1802641720, 1980128},{0, 67108864, 0, 1110804928, 933576812, 1422629, -384594996, 2, 71846912, -1961983063, 8, 1114112},{0, 50331664, 0, 1076527104, -145036924, 760980, 1880956216, -1073741821, -1965398107, 2140391604, 6, 546816},{-2147483648, 1, 0, 738197504, 1091433732, 551005, 886260280, -1572601842, 773907, 0, -1036255232, 1781152},{-2147483648, 1, 0, -1342177280, 1363517701, 1000361, -1811939328, -472897711, 1943413, 2100318660, -2147483637, 1773893},{0, 65, 0, 335544320, -1849124687, 1353808, 1610612736, 1610612740, 1174543230, -1495284684, 26, 849920},{65536, 48, 0, 1375731712, 824279051, -1014061531, 1444479372, 1074003988, 1384379, -438353920, 27, 1974272},{268288, 83886112, 24576, -1342177280, 1547482233, 868444, -1027967064, -2147483625, 1774515, 461365248, -1750335484, 269264},{69632, 48, 0, -268435456, 475447309, 1015910937, -2032065816, 1447297038, 1341354, -1538549892, 1467744282, 221213},{0, 33554480, 4096, 1879048192, 1812551692, 549473797, -1569711135, -1684013027, 551186193, -617918183, -605478697, 1976963},{196608, 0, 0, 1140850688, -660422214, 693144, 1134188440, 14, 44032, 899842048, -2129133542, 1165202},{-2147221504, 33, 0, 1880522752, 624603410, 1649368557, 1807646064, 592196609, 1217272739, 1297177300, 1523843735, 1466705},{6144, 0, 0, -1342177280, -1862137315, -1244878758, 394310112, 1264362241, 381020, -469762048, 1184366605, 535838},{0, 50331648, 128, 405471232, -148443902, 1876122772, 2027887153, 14, 1901735936, 1451117717, -1183580156, 1527722},{0, 16, 0, 100663296, -1530781086, 638754284, 491394185, 1392070350, 1374105, 1632550912, 1073741836, 1780646},{-2147483648, 33554433, 0, -1442840576, -1420713725, 1031712, -1321120276, -397127206, -523373661, 1116968048, -1804548274, 950698},{268288, 32, 0, 0, 715530659, 1963834605, 1942253904, 1525415950, 1373096, 1891027624, 1327019649, 1165596},{0, 32, 12288, 1075380224, 1462137923, 2119588821, -304261243, 382041693, 1781705, -239150228, 395074267, 569908},{0, 16, 0, 101220352, -1537547629, -942967982, 753028640, 1311040023, 1542748, -1610612736, -2147483636, 733348},{2048, 50331680, 0, 1754300416, -1143321940, 1988981542, 171175588, 305659934, 1151017942, 400196361, 1528369563, 1329586},{0, 50331680, 0, 1342177280, 2068979970, 1074947431, 775405580, 11, -1433687488, 937347900, 188235806, 1930296},{0, 0, 0, -1037631488, 666248117, 386554449, -964354648, -2147483631, 239663, 31113588, -1049624559, 774617},{196608, 16777216, 8192, 0, -145307286, -1265541676, 1183518077, -2112085615, 566425827, -1908961732, -1073741804, 920540},{137216, 67108864, 0, 1342570496, -1488838371, -1982444690, 985461188, -2006712303, 1498935434, -2095330288, -954728447, 1565811},{137216, 0, 0, 34242560, 960941676, 667532831, 1675256784, 500695066, 1247506, 1494359512, -1073741804, 967114},{131072, 16777216, 384, -1409286144, 681701483, 327767599, 1188024645, 1566572546, 634256867, 855933784, -479861861, 932387},{0, 1, 12288, 402653184, -1998921444, 936266906, -438270308, 1910767643, 1165233, -1726069868, -2121006820, 1334205},{131072, 67633200, 0, 1073741824, -178407803, 2081526492, 1675255101, -575026940, -909876261, -1572602355, 11, 1969152},{196608, 64, 0, 2424832, 1766924715, 1406622619, -1977739311, -1669857266, 903727, 1642102784, 1577582595, 249213},{0, 50331664, 0, -1006632960, -145309683, 1838324816, 91592533, -786694137, 2052578080, 722570928, 30, 460011},{0, 16, 16384, 1174405120, 1957831237, 1854575469, 738919552, -2037383143, 1746850, 2115076096, -1073741801, 1850957},{-2147483648, 33, 4096, 604536832, 2055903338, 621485, 0, -145995584, 1120995, 1677721600, -726138858, 1829474},{0, 68681808, 8192, -1342177280, 1453775036, 1196531781, -193538939, 1716054932, 1564772259, -1753160036, -1901518650, 72527},{0, 17874944, 16384, 805306368, -1677297583, 222340, -736394916, 1285124433, -406630782, -682526898, 1373139546, 403167},{0, 48, 4096, -1339588608, 1506953483, -489202283, 1604721028, 1528148235, 911056, -1926149216, 20, 1172992},{71680, 0, 0, -1844871168, -1254219236, -1323977176, 853486713, -2085878566, 1746140, 339247104, 27, 320735},{0, 0, 0, 1107296256, 1633559395, 1275051, 1545404416, -1849384117, 1371884, 1409286144, 17, 1159168},{0, 16777264, 0, -2147483648, 373359181, 892079, 1641955328, -1640759267, -754021532, 1937235513, -2147483628, 1961438},{0, 0, 12288, 1879048192, -2133696483, 821412, -195772416, -1073741819, 1372494, 816104780, 308827339, 1766259},{65536, 0, 0, 1140850688, -190676116, 1221546, -429154788, -775301609, 486691, -216228324, 27, 960512},{2048, 0, 12288, 1476395008, -1473871333, 941410, 652359684, -1073741810, 2145078357, 950787585, 1075175435, 733760},{0, 16777248, 0, 1879048192, 1495401228, 957851, -1467301888, -1897136125, 1318955568, 1250399477, 1213762388, 1779223},{-2147483648, 65, 8192, -1332740096, 120693010, 567250327, 48368768, -478662524, 1226718, -1454389668, -1795424245, 230024},{0, 0, 12288, -1340833792, -707648998, -766536790, -1591943655, -568852475, -2028876692, -1350678368, 29, 774656},{-2147483648, 64, 0, -2056224768, -1672846419, 684888, -807567360, -39321571, 1930785, -1311211520, -1899636004, 250920},{196608, 0, 0, -1040187392, 448168563, 290635169, -958407115, -2107375599, 853045, 0, 1073741824, 476119},{-2147483648, 50331648, 0, 704643072, -1861920765, 1206992, 1610681232, 536870941, 1956626, 1541521408, 111411220, 1828920},{131072, 0, 0, -268435456, 551100437, 1409251, 1205436416, 17, 125952, -268435456, 1517821697, 1744302},{262144, 16, 0, 807665664, 1342527665, 893139, 1458134548, -569114616, 2136074032, -850979752, -1660682237, 126185},{0, 16777216, 16652, -1342177280, 1275246666, 754448, 205462200, -1793563772, 1268629265, 257000464, -1210158946, 1739738},{0, 32, 16512, 100663296, -189125278, 1201578, 832061440, 1073741850, 221768, 174671068, 1622699742, 213885},{65536, 1048576, 0, -973078528, 1463186058, -1307148759, 1541414349, -618575017, -1252130340, -1290666547, 473694222, 1793501},{0, 16777216, 16384, 1140850688, -1406295180, 1353730, 1297040968, 6, 960803, 457676024, -1073741823, 200311},{0, 17874944, 0, -503316480, -1530849933, 1220076, 1476395008, -875526770, -1122546034, 531494074, -1049624555, 771099},{262144, 0, 8576, -1677721600, 1278615725, 1067077, 54607872, 300417041, 875850, 1704628712, -298292454, 1375006},{0, 67108864, 4364, -2147483648, 1277311050, 1023109, 2108184408, -1073741811, 919924, -1237723544, -1376379576, 1170152},{0, 0, 0, 1174405120, -794164595, 941208, -1006632960, 1073741841, 836441877, -793343300, 1073741838, 1765405},{131072, 16777216, 0, 1879048192, 1102405653, 1144225, -1284661708, 26, -560122880, 400481653, 27, 1542144},{0, 50331648, 0, -266731520, -517916645, 1138714, 353370112, -623378405, -1383729068, -210560231, 1430538714, 1563005},{0, 67108864, 4096, 503316480, 1373224972, 880785, 1073741824, -1669595116, 960631, -1746894848, 1, 1960556},{0, 50331664, 0, 67665920, -1185763732, 610846, 967937648, 346554379, 1373109, 867254272, 11, 712704},{-2147483648, 17, 0, 805306368, 537212957, 1083547, -1140850688, 682640068, 1121045319, -2000823620, -1698938552, 777355},{262144, 16777216, 12288, 805306368, -2130298735, 189642088, 260075044, 351620882, 190119014, 46813856, 1073741854, 242187},{0, 0, 8576, 33554432, -1767207277, 1006800, -805306368, 141819910, 1565834, -161824768, 1909555348, 241342},{69632, 0, 0, 1610612736, -380001532, 1002982, -1439189252, -2026373109, 1921400, -29538500, -2025848812, 168410},{262208, 0, 0, 805306368, 562465369, 659581091, -673074738, -1794899963, 875936, 760233984, -617799141, 919605},{137216, 67108864, 0, -1342177280, -2136604531, 470717082, 601734036, -1684785391, -1180820479, 467092353, 23, 228352},{0, 48, 8192, -1040187392, -1188954035, -989164774, -236872407, 354269505, 1737574943, -1652583140, -670280422, 1981409},{0, 35127296, 0, 1107296256, 667000948, 1292845, -643022848, -988282851, -884748834, -222730247, -2147483631, 150956},{131072, 0, 12288, -1844034540, -113939795, 295149084, -1085176259, -1699904931, -1429991314, -227339795, -1073741823, 1764126},{0, 33554432, 4096, -1342177280, -121568501, 1413736, 372529876, -1073741794, 1676365, 1912898708, 1150563476, 957347},{0, 524320, 0, 1191215104, 957011387, 625567, -1071069652, 82600730, 739580844, -1035912360, 26, 180323},{65536, 32, 0, -2046820352, -710541174, 1472042, 652907020, 105644033, 454264, 2013265920, -2147483642, 1341775},{4096, 48, 16384, -2113929216, 1472615451, 428455121, 601892956, 27, 1953314, 538690108, -1073741822, 263715},{0, 67108864, 4096, -2046820352, -870137268, 1411074, -1189178112, 301727769, 1729872, 1994622644, -1073741823, 1376982},{262144, 16777217, 0, 469762048, 1219945289, 46616, 531301592, -1399062526, 774844, -1951507748, -1762809714, 914805},{196608, 0, 0, -1442840576, 1085612547, 1152417, -1558880768, -2147483628, 1174198, 766451204, -614465521, 708657},{0, 32, 12288, -268435456, 547700906, 1263448913, 954764913, -1691766243, 241630, -1998028800, -1073741801, 1750894},{196608, 0, 0, 1140850688, -1069219478, 1463210, -206733312, -953155558, 1930899643, 206179260, 1073741830, 558195},{0, 68206592, 0, 570425344, 1789993245, 1293467, -294104024, -1073741795, 1191635002, -337396245, 38535195, 961594},{0, 33554448, 0, 1778384896, -188644597, 1116619876, -1588623792, -2077229050, 1780144975, 447941200, 67371035, 1563242},{65536, 32, 0, -2046820352, 1342838909, 611409, 512425984, -1073741794, 1168299, 430702592, -624144828, 312459},{0, 0, 8576, -2113929216, 1790784619, 1716999331, 450499836, -1853358053, 46513, -172912248, -297946540, 1967946},{0, 17825792, 0, 809140224, -2004535293, -661824892, -463779679, 23, 486813184, -542381959, -1008467957, 448984},{0, 48, 0, -334102016, -391470563, 889562, -1981856792, 1195237207, 1473576509, -1713711335, -2147483646, 1564029},{0, 48, 8192, 503316480, 1348059410, 1528425, 78907592, 21, 576195252, 137741009, -1073741810, 1168086},{0, 0, 8192, -2033122752, -196771421, 1291602, 473374236, 0, 1921220608, 231346648, 1536761246, 1945117},{0, 16, 0, -402653184, -1858747637, 1049736536, 360711584, -617349090, 1378264, 802741704, 27, 1903071},{0, 0, 8192, 1075118080, -616397910, 752536, -872415232, 3, 528384, 1551958016, 2, 1974913},{0, 16, 16384, -2080374784, 617677741, 900189, 1011843072, 26, 2044009984, 1460782917, -968514532, 1166161},{0, 50331664, 0, 1879048192, 202225690, 2069127303, -651735412, 233621207, 2099113697, -1683793495, 14, 1755881},{266240, 16, 0, 805306368, -1531591815, 1058319044, 1330757116, 401080325, 1117433423, -295494112, -975699951, 1786946},{196608, 0, 4096, -2080374784, 952022123, 1489509, -541097984, -1678162876, 1146806087, -1994171499, -771489785, 215786},{131072, 16777216, 12288, 1879474176, 1960381972, -2104338913, -1037959035, 447564378, 289883563, -1022062308, 1417224450, 1954321},{0, 18350080, 0, 1140850688, -1448771445, 1209694, 1677721600, -771734182, 386808023, 55556556, 21, 283648},{-2147352576, 50331648, 0, -1622114304, 2025459021, 679141, -1082549448, 987620225, -1299457502, 1064670973, -1641545726, 320946},{6144, 0, 0, -1342177280, -524148220, -1232569112, 52342588, 21, 954368, -1870921728, 503694286, 1136814},{0, 16777264, 0, 0, 1471529618, 701651, 566214656, -1752609317, 832222952, 258986977, 465567758, 1302976},{0, 48, 0, -1073741824, 1625104978, 814097, 812843008, 1073741847, 1765962, -1131921408, -1037295029, 397741},{0, 48, 0, -1072136192, -146169180, 1397328, -115441664, -2147483646, -1059198406, -328499195, 17, 1838519},{-2147084288, 66, 0, -1810202624, 347191385, 1700020359, -206724052, 733899265, 1744415, -122617856, 185633866, 736322},{131072, 18350080, 0, 0, -1747604339, -740912240, -743711255, -1645740015, 334989, -1354275640, 14, 1755136},{65536, 64, 0, -265715712, -1042735091, 678736, -100663296, -636747756, 1552159354, -1918838944, -990546418, 1159400},{137216, 16, 0, 1879048192, -358481900, 517127554, -566024775, -957087733, 1752862, -1457699076, -1848377336, 1566782},{196608, 33554448, 0, 0, -1456607734, 1040812826, -29539347, 142344212, 1776170, 1060309972, 14, 775168},{0, 50331648, 0, 1881538560, 732086530, 684899, -528515072, -769073651, 919767, -771751936, 49107089, 1936950},{0, 0, 4480, -1342177280, -598334971, 310940590, -164101516, -2138308579, 1973266, 1946157056, 539350851, 1564537},{6144, 0, 0, -1778384896, 279265820, 487828769, 1129347897, 11, 1951872, -1390604780, -837550075, 1573997},{0, 0, 0, -2046820352, -1589550747, 1152490, -60391288, 20, 156672, -615513976, -1064828911, 250084},{0, 0, 8192, -2113929216, -1683913851, 691098, -729235456, 62700875, 131960548, 538084296, -1054341106, 1973959},{196608, 16777216, 8192, 1879048192, 1453457426, 2072925609, -1617195540, -1073741810, 1717435, -1563997248, -930611186, 959357},{-2147483648, 33, 128, -637534208, -147771054, 1289508, -1744830464, -32485225, 1122169, 0, -52069952, 1721169},{131072, 0, 0, -258932736, 1373217029, 496063393, -616065979, 23, 495397888, -1388031483, 306708494, 955001},{0, 0, 4480, -268435456, 1006802946, 1200263, 565362688, 17, 1905992704, -218967175, 1956120791, 274348},{0, 16, 16384, -1409286144, -1856683157, 1017304, -98762752, -2147483621, 1328929, 0, -1713627840, 571302},{-2147155968, 50331712, 0, -268435456, -785792998, -376406680, -1217313964, 928629760, -2116749397, 400720740, -1073741823, 151785},{131072, 0, 12288, -268435456, 469940226, 610375, 988348416, 1204113870, 284404, 1487896576, -719559535, 1377974},{0, 67682304, 20480, -1073741824, -2025151892, 1538668, -1989065680, 1073741847, 545526084, -1347241241, 1143818077, 476092},{0, 50331648, 0, -1442840576, 279290372, 679129, 683655168, -1950564395, -1072786913, 102910088, 30, 1520640},{0, 67633200, 0, 1879048192, 189964802, 1145557, -1473209260, 1536950275, -1155847227, -1690420364, 1269861915, 1835520},{0, 0, 4096, -2080374784, 1077289875, 1416145, 1170538496, 1521605403, 724395, -1313259520, 1549008925, 1761158},{0, 17825792, 0, -1341882368, -1210932469, 1152404, 876707840, 4, -1211878400, 253682892, 28, 752640},{0, 524320, 12288, 805306368, 1237922060, 1658153625, -1334127396, -995622905, 275176, 313785060, -623116277, 1380072},{2048, 48, 0, -268435456, -519235557, 1092866, -341056532, -1651769315, 778863, -395313152, 23, 376832},{-2147483648, 1048640, 12288, -268435456, 1277604277, 693121, -268435456, -492271615, 835072928, -1888078879, -2074607602, 1779261},{65536, 0, 0, -2046820352, 469874837, -2041823101, -298875151, 140509201, 517481658, -701099535, -1073741807, 1599674},{262144, 0, 12288, 805306368, -259884971, 1179226268, 570572944, 2, 288768, -700022784, 1131949771, 1964600},{2048, 0, 12288, 1140850688, 71224941, 1532072559, -488589308, 461111309, 1851841, 364969984, 471186076, 1379293},{4096, 0, 0, -1342177280, 1353278213, -2113029101, 736227029, -1791492095, 1401056264, -789751775, 356253699, 972162},{65536, 0, 0, 100663296, -1235557812, 889940, -767835812, 17, 927744, 382566532, 1073741838, 776329},{262144, 16777264, 0, 67665920, -1681266076, -1085454948, -1952230867, 1073741838, 959423, 60611432, -720547691, 913607},{0, 50331648, 16384, -1342177280, 1619077147, 1075371, -676901828, -1073741813, 1851587, 736119804, -2147483647, 472999},{0, 48, 0, 1140850688, 1700110658, 1863415255, -1390112304, -733741042, 956025, -1040187392, -2147483637, 1342752},{264320, 50331648, 0, 1879048192, 440330, 1406236059, -1548961805, 6, 1350972, -149793408, -1751295977, 997810},{0, 0, 0, 1174405120, 1364910226, 1345617, -1275068416, 20, 1356800, 1744830464, -1073741798, 1700913},{0, 50331648, 0, -2147483648, -2134760886, 768922, 417890304, 454295579, 1898626, 639979164, -2147483647, 1979445},{65536, 33554496, 0, 1174405120, 201758738, 802819, 175936096, -1962147819, 568085, 1593103012, 1073741828, 955690},{131072, 0, 0, 1543503872, 27631876, -95245039, 1525782372, 249123607, 274742, 1694269440, -680985452, 958193},{196608, 33554432, 0, -1342177280, -795957228, 571061154, -1823292888, 14, 1624579584, 1869827009, 1443717131, 786571},{0, 50331648, 8192, 1075314688, 618293860, 768875, 1677721600, 1073741833, 766102, 109992936, -1021537700, 1543738},{0, 0, 0, -1006370816, 1354310581, 678875, 70664208, -964599722, 1744209, 626901872, 21, 1750016},{6144, 16777216, 0, -1342177280, -1593462757, 986799378, 1472311416, -1012924388, 1068295, -1291337132, -799277045, 270599},{0, 16, 384, 67108864, -632927164, 1422246, 1006632960, 129096715, -1935822237, -1914959088, 887111246, 1857204},{4096, 48, 16512, 805306368, 78991618, 1209837, 918429696, -1853358076, 780158, -652705792, -536870907, 1564588},{0, 524288, 0, -2080374784, -1180032156, 949530, -939524096, -2147483629, 776330, -420912168, -1073741798, 184636},{196608, 32, 4096, -1342177280, -603604972, 1138692, -1900406744, 140771357, 1169974, 0, -778567680, 1176113},{131072, 0, 4480, 1879048192, 1275410564, 273563651, -634420120, -1073741813, 1834425, -2076730372, -532938749, 1304133},{0, 33554432, 4096, -1342177280, 537319442, 1132779, -239009792, 28, -1159981640, -228745759, -2147483631, 1600384},{0, 50331648, 0, -245366784, -1598643683, 298748952, 1968410904, 404811074, 2110024253, 988417684, 18878081, 1121395},{0, 16777216, 0, 1778384896, 1099296772, 616605, 700792832, -610271218, -1986260275, 370559960, -2147483620, 246213},{0, 0, -1744830464, 103450176, -1805817203, 949100, 0, -1687420928, 426207, 13451264, -1073741803, 1718685},{0, 48, 8192, -603979776, 270639379, 1413737, 296246088, -1649410018, 80847, -1275068416, -628621283, 777132},{0, 67108864, 0, -1342177280, 12952324, 542873, -159186100, -765983525, 501063, 109248512, 55050240, 962691},{0, 0, 0, -2046820352, 279355978, 1225513, 1065096348, 12, 1008640, 671088640, -716963813, 1124668},{137216, 0, 0, -2113929216, 992084108, 147672405, -616269304, 17, -1149202432, 1546771481, -2147483644, 37313},{0, 0, 0, -1342177280, 1373184514, 557145, 1275068416, -1026026798, 161304629, -2082253748, 21, 1330176},{-2147352576, 16777217, 0, 1879048192, -150808477, 572434, 253073164, -278646443, 1731141, 238081792, -972029931, 1206275},{0, 50331648, 0, -2080374784, -63569524, 566182, 436207616, 1336760731, 1294675, -1620230144, -2147483634, 1338732},{0, 0, 8576, 805306368, -1420410622, 871644, 805306368, 19926081, 928462169, -1486863492, 578289682, 956087},{0, 0, 4352, -1342177280, 25835524, 629585, -1342177280, -2147483637, 209038, -902117080, -1589379057, 991094},{0, 32, 12288, 1879048192, 977412355, 1004453, -1917744984, -706691711, 770614, 262881280, 1372110422, 143282},{262144, 32, 12288, 805306368, 436328529, 884805, -1969852320, 0, 766525, -519749632, -2082461822, 1842746},{65536, 33554432, 0, -1338605568, -1530494964, 1290986, 112869376, 1215823894, 1045085660, 649305536, -2147483627, 256187},{196608, 32, 4096, 1879048192, -1073031157, 1137298, 991515096, 4, 1080832, -268435456, -974579311, 1081214},{-2147483648, 33554449, 0, -503316480, 333939, 1413723, -381842472, -472302206, 1950440, -503316480, 20, 570368},{0, 0, 0, -973078528, 1364894130, 610329, 1638350848, -1691615229, 209176, -1534649556, 11, 1175552},{0, 16777216, 0, 100663296, 1359378610, 1220611, -2077196016, 20447235, 227770, -435929088, 19, 0},{0, 0, 8192, 1174405120, 3252548, 961705, 360742912, -1682857764, 1958351, -134217728, -633602044, 1601401},{0, 0, 0, -2046820352, 1359100053, 1337441, -797130752, 3, 1834564, 537837568, 1073741825, 164073},{196608, 32, 0, 1879048192, 277501098, 1270433, 303467508, -976486372, 1981552504, 953598913, 205258766, 1576644},{262144, 0, 4352, 805306368, 1342811273, 1327315, 850840384, 4, 537003008, 954240364, 972328218, 1121810},{0, 68681728, 0, -1845493760, -793075115, 1021016, 134217728, -603343332, 1921449, 45981696, -600047604, 1858529},{0, 50331648, 4096, -2080374784, -63881109, 1465696, 2085765120, 440401940, 1225859, 183179840, -1018421924, 1379962},{0, 1048576, 0, 1174405120, 8476692, 1219859, -669826860, 19, 1975596032, -1213402995, 389634525, 1130826},{0, 0, 0, -1039630336, -1856896174, 961690, 469762048, 1073741848, 286086, -1140254620, -633319397, 213414},{65536, 50331648, 0, 67108864, 1788985421, 621435873, 803423069, 27, 1930240, -2043805696, -1073741803, 77833},{0, 17825792, 0, 101089280, 1216714882, 678493, 3201548, 23, 1415168, 463921220, -636464612, 1137910},{65536, 0, 0, -268435456, -779802619, 1409196, 794771456, 1, -499122176, 1330042573, -566493164, 1297887},{0, 50331648, 0, -2147483648, -1856896597, 1464976, -938377216, 1121452032, 1415223, -1442840576, 1092357074, 1521683},{262144, 35127296, 0, 335544320, 1344575609, 868445, 1800292596, 4, -1269020672, 1794964136, 23, 738304},{65536, 0, 12288, 301989888, 21381133, 1399441, 842451728, 1073741825, -1010102081, -1799518052, 205258753, 1446543},{-2147143612, 1, 16384, 805306368, 1816180849, -1767328790, 585984946, 1657880344, 1057205780, -1473330215, -799510141, 1392436},{0, 50331648, 4096, -2147483648, 399868523, 1068437, 948600832, 11, 1145809372, 313394152, 22, 1779200},{196608, 32, 0, -2147483648, -1716412044, 679454, -2107714912, 16, 1082154, -325695204, 1381761047, 1159318},{131072, 0, 0, -268435456, 1346749203, 508848225, -1036151827, 1529433949, 194878, 1080606720, 299892755, 1779007},{0, 16, 8192, 100663296, -1422745582, 619362, -798932992, 1215623566, 1176250, 404504700, -1794106161, 1171281},{0, 48, 0, 2655776, -995986772, 683500, 2021670912, -2128867901, 777732, 484707860, -1073741823, 231473},{0, 0, 4480, -2080374784, -441281652, 285911642, -397934300, 411151645, 1781717, 603979776, 2048503169, 223007},{0, 32, 12288, 1107296256, 958537890, 961369, 1088290816, 1092620036, 1836777, -2004988400, 1207959554, 81469},{137216, 0, 0, -2147483648, 1439834452, 834983, 394321920, 205307868, 931900, 0, 394882496, 884759},{0, 33554432, 0, -465960960, -1069178604, 1397650, 159335748, -671350758, 919723, 582386184, 1, 884736},{0, 0, 0, -973078528, -1859559276, 1065058, 1709050812, 1523437787, 1973719, -1744830464, 8, 1959100},{0, 32, 0, 806813696, -2118770667, 1422496, 268435456, 314423388, 1719019, -582483124, -1073741817, 204225},{0, 65, 0, 809041920, 876749061, 1466987, 192233688, 1610612764, 1083881435, 1091163297, 17, 1498112},{0, 0, 0, 100663296, -1061797262, 1350242, -1983882248, -1684537320, 1721252, 1476395008, 1073741852, 1582533},{65536, 0, 0, -1342177280, -237699059, 813212, 921600000, 1, -288430080, -2010201808, 10485789, 1980470},{196608, 17, 0, 805306368, 717651978, 627501, 1593249304, -1605805244, 1599425, 1567637504, -873463791, 200929},{0, 48, 8192, -1677721600, -1071275758, -1319795760, -666427872, -691150253, 1331014, 0, -887582464, 78687},{0, 0, 0, -1006632960, 1352811372, 1462873, 1946157056, 1073741827, 1522011, -535609344, 12582914, 1708557},{0, 0, 0, 1177223168, 1078534557, 1530531, 1169063948, -1706819558, -2120740642, 350129129, -1073741798, 1709486},{0, 0, 384, -1342177280, -1056101118, -1856993176, -1732408328, 1, 739328, -1263239168, 1668284424, 73235},{131072, 48, 4096, -402653184, 104190355, 1421905, 1241513984, -2082996196, 1952098874, 1177473112, -749731829, 1370671},{0, 16777216, 0, -1342177280, 1096123149, -607273963, 314219969, 1572193291, 718916, 1049313280, 12, 736256},{0, 16, 0, -1073741824, -779790221, 1132708, 0, -920649720, 1307518, 1629339648, -1911291886, 390369},{0, 50331648, 0, 1140850688, -794689356, 1220074, -1006632960, 36445908, 1354958953, -954334675, -1073741795, 253264},{264192, 0, 0, -1338605568, 1149605892, 366035093, 858401700, 8, 134333440, 1720161552, -1054343159, 400402},{0, 32, 4096, 1073741824, 958530412, 631773, 939524096, 227616142, 1780238, -2012949492, 1073741827, 1307457},{0, 65, 0, -771751936, 1891172435, 1468641, -1476395008, -1116363945, -1296002319, -310322383, -629669859, 1686912},{0, 16, 12288, -2147483648, -788121436, 957016, 162709504, 1301394062, 73346, -735506788, -1073741821, 229245},{0, 0, 4096, 100663296, -1489878374, 1007264606, 652447120, 1, -1010042880, 1970837228, 1, 1759744},{0, 48, 0, -2147483648, -793107804, 1264984, 148439040, -2147483634, 74422, -799916032, -636485622, 1570900},{0, 0, 0, 100663296, -1061830020, 1280684078, 500243153, 1073741854, 296274, -1981917916, 29, 1759232},{0, 0, 0, 1174405120, -1054793645, 1353826, -1312735232, -1020150962, 1343540, -469762048, 7, 1230848},{0, 48, 128, 1509949440, 72450573, 965741, -2080374784, 346140250, 1842964, -1318135068, 1947825552, 771038},{0, 0, 0, -1073741824, -2126101588, 1335392, 603979776, 15990785, 1729554, 96370688, 475529244, 1686974},{0, 0, 12288, 1140850688, -1068940965, 959714, -1725906944, 1073741853, 562809121, 943065245, -823346146, 80431},{0, 48, 0, 1073741824, -2127486637, 1152288, 0, -687514688, 1601301, 2016477260, 15, 783360},{262144, 85458944, 0, 1141178368, 1471316330, 750627, -414787892, 19, 1610677248, -367840247, -1053294573, 594963},{0, 0, 0, 805306368, 833995266, 1138789, 947964108, 1221853207, 1424512, -327106560, -1999110142, 925239},{0, 0, 384, 805306368, -522591742, 688746, -402653184, 26, 1577984, 482263040, -535822312, 728035},{0, 33554432, 12288, 33554432, 1699872843, 888165, -527335424, 1073741835, 757853, 915244492, 1221090625, 75405},{196608, 16777248, 16384, -1342177280, -603580254, 1057187332, 1178239960, -2111561766, 911906, 373343236, -485740582, 280494},{0, 18350080, 0, 1879048192, -388890107, 1477006166, -1316579283, -664272885, -1328854386, 1925475132, -2147483645, 1410388},{-2147352576, 65, 0, -503316480, -1604755052, 965482, -215072768, -1476115565, 1052904197, 340821049, -2077933874, 328783},{262144, 48, 0, 1107296256, -1808145756, 882029934, -807669084, 197432026, 1951518, -1799601344, -1071382522, 1222950},{131072, 50331648, 0, -2113929216, -1448169628, 543580, -1440989184, 18, 311948113, 1854424608, 8650761, 763927},{0, 1048592, 0, 100663296, 962144395, 939483, -796606464, -1908622133, -595448264, 238936144, 121634837, 1135893},{0, 0, 0, -2046820352, -514514566, 550946, -268435456, -627310573, 1961394, -1986145468, 29, 1718591},{131072, 0, 0, -973078528, -1538932333, 143895826, 595531688, -1745874559, 250921, 335544320, -844890111, 1316576},{0, 0, 0, -2113929216, -1054760052, 619808, 2026094592, -1073741823, 1542511, 249187328, 1073741848, 932924},{0, 33554432, 16384, -2046820352, 1791107402, -1551057691, 783713613, 1073741851, 2140409131, -1562752287, -736886770, 1976032},{0, 0, 0, -2046820352, 1086464683, 550931, -1744830464, -1993605091, 1959062, -733427352, -2147483622, 1974737},{0, 0, 0, -2076475392, -799686275, -2066707822, -381154436, 1073741831, 1841336, -872415232, 18, 964030},{0, 50331648, 0, 1610612736, 1093771546, 955473, 1095375860, 1412001745, 1386252, -411722900, 29, 1833984},{131072, 0, 0, 1174405120, 1079345538, 1490001, 1309802496, -1073741821, 1836047, -574710796, 25, 1730560},{0, 0, 0, -973078528, 282477164, 1471017, 357351424, 505498770, -505747914, 482085045, -1073741821, 1926241},{0, 50331712, 0, -1342177280, -782884837, 548960, 1571340288, 445138897, 1641143857, 1511413513, 28, 1015808},{0, 32, 0, -2145779712, -1698331797, 1000614, -1336654348, -685411945, 1981306, 0, -1764663232, 1339713},{0, 50331648, 0, -1040187392, -2142920077, 1219944, -722616320, -633864184, 931663267, 527685080, -819924530, 196000},{0, 50331648, 0, -1006632960, 1763778898, 1389473063, 272733933, -630718464, 1852838, 465852152, -636747765, 81838},{0, 0, 0, 102367744, 1429586554, -1009628073, -719729600, 246764936, 1456576704, -731330543, 5, 1403904},{65536, 32, 0, 100663296, 1482354253, 1201243, -349487104, -1804254003, 1709600, 472023040, -1008979773, 1722938},{196608, 0, 8192, 1779827328, -333287549, -619213404, 1264127504, -1790181365, 1451965782, 829853197, -1062897407, 779795},{0, 0, 0, 1174405120, -1062641044, 1876143250, 82057053, 5, 922624, 249681752, -867172348, 536878},{0, 0, 4480, -1842872320, 2067681634, 895709, 1778535240, 24, -1224523776, 1085376888, -1310430773, 1410747},{0, 33554448, 0, 1879703552, 2067858194, 873821, 269008896, -2147483627, 390347282, -289765240, 1073741843, 116834},{0, 16, 8192, 1073741824, -408329339, 881452, -2000896000, 3, 1317783040, 1427441477, 1312817152, 1223301},{0, 0, 0, 1174405120, -246341235, 1032679440, -304506067, 29, 1750016, 966738956, 26, 265216},{0, 67108864, 0, 808779776, -522903431, 181690522, -735444716, 3, 920576, -287534424, 14, 1222951},{0, 0, 0, -253493248, -782630139, 1353816, -210206720, 1227882515, -1131564868, 1010581888, 14, 1513472},{65536, 0, 0, -1073741824, 1363256245, 543657, -209742836, -2058015785, 897199, 201326592, 14, 748544},{0, 0, 12288, 67108864, 3522986, 1624347609, 957649185, -704291388, 276722, -2080374784, -1786424107, 803394},{0, 0, 0, -1073741824, 290866100, 819281, 1409286144, -1073741807, 520434, -1256734720, 192972110, 1344813},{-2147483648, 16777217, 8192, -301989888, -1235602028, 1068308, 0, 1950446976, -1190564898, 588094457, 1420128670, 1760020},{0, 0, 12288, -1073741824, 10560082, 1346393, 92706864, 1, 0, 1772044288, 1546225370, 1842706},{0, 0, 0, -1073741824, 558719859, -683055019, 1613960393, 3, 1973248, 549060608, 6, 0},{65536, 48, 0, -1342177280, -802782694, 1422040, 103874920, -1761072740, 1858297, -936640512, 2, 1139042},{0, 48, 0, 1879048192, -1060970469, 1353900, 829527980, -1764728938, 772930, 1879048192, 20, 347136},{0, 0, 0, -2080374784, 281617325, 891665, -1891118412, -1015439014, 1523037, 2013265920, -2147483624, 200010},{0, 0, 0, 0, 1104568754, 821413, 1543503872, 1, 1503577, 2041495552, 24, 1722434},{0, 0, 4096, 0, 289997723, 1421921, -1722431128, -915893487, 430422, 0, -1073741824, 991972},{0, 16, 0, 1879048192, -1070169334, 1209043088, 833149576, 3, 1193035264, -1405238499, 3, 1321984},{0, 17825792, 0, 1879048192, 25866506, 1220009, 1121883472, 12, 1925185536, -1151934155, 395051022, 54469},{0, 67108912, 0, 0, 1085653626, -53035687, -1327413200, -1882916467, 142197, 1064406588, 26, 0},{0, 32, 0, -1342177280, -1867915243, -1282522902, -1607185560, 1078504966, 1403678, 0, 0, 0},{0, 48, 0, -2080374784, -793083731, 1220066, 2014478336, -2002253567, 1308346, -939524096, -2147483647, 1381474},{0, 0, 0, -1073741824, 567959996, 1155243, 1552238408, 0, 1134592, 536870912, 21, 232637},{0, 0, 0, -973078528, -1858960980, 1150992, 2030359624, -1807220720, 1718688, -1071017408, 46729282, 1308083},{0, 67108912, 0, 805306368, 1363329377, 565267, -1461662244, 2, 1370624, 461707316, -2135587566, 251921},{0, 0, 0, 1110706464, 1439291012, 813737, -1921875968, -2084246719, 933084, 0, -1073741824, 1962872},{0, 0, 0, -2046820352, 1087816266, 750417, 0, -2057830400, 920796, -1430861044, 315097106, 1572161},{327680, 0, 16384, 1879048192, 1093051289, -1160738715, 257969116, 8, 1107968, -883027644, 11, 580096},{0, 0, 0, -2046820352, -526237110, 1083418, 1427587072, 283639816, 963713, -2068316160, 20, 1239040},{0, 84410432, 0, 1879048192, 22591673, -1797953315, 997562152, -1684799484, 243652543, -614960827, 1073741832, 610451},{0, 0, 0, -2147483648, -2127133780, 1083480, 0, -1673522624, 1730976, -536870912, 26, 1754112},{262144, 16, 0, -2046820352, -262749556, 1526300, 1050017792, -764411893, 1353512, -920076288, 505534923, 222260},{196608, 67108864, 0, 808026112, 741382209, 1083463, 1512701952, 28, 1679232044, 185995169, 1097859077, 1601073},{65536, 0, 0, 1174405120, -1876336027, 889936, -814938804, 388057684, 1339716, 962434212, 22, 1552384},{0, 0, 0, 1073741824, -1581129075, -2062716846, 1010276921, 23, -2079023104, -533605351, 21, 1594368},{0, 67108864, 0, 1161232384, -1063074925, 1083434, 1766637604, -1021038118, 1422766, 1107296256, 348938830, 1504279},{0, 67108864, 0, -2143617024, -1059741053, 1538600, 1824686080, 21, -292804608, 241782532, 1276702788, 1154390},{0, 0, 12288, 1142554624, -1163788150, 1291412, 805306368, -997898493, 240701, 0, 445465664, 1854004},{6144, 32, 0, 1744830464, -148791022, 328226134, 1793830412, -786623351, 1934978855, -512175472, 287077197, 1405225},{0, 0, 0, -973078528, 1093288090, -1794095005, -915042364, 13, 933013, 754581504, 23, 606208},{0, 0, -1207959552, 36964768, -1188680013, 687316, 217071616, 11, -281018368, 1286851436, -2147483648, 215280},{0, 0, 12288, 1073741824, 1096122803, 1132001, -1469939712, 1073741835, 117214, -2125373968, 1562116097, 924299},{0, 0, 0, 67108864, -1061780619, -610960816, -435809967, -1073741807, 774277, -1938481920, 3, 1949696},{0, 0, 12288, 1107296256, -1874754963, 1135528, -1046249472, -1861676990, 1070122, -1110769664, -952775716, 77575},{196608, 0, 0, 1107296256, 1348051588, 1536537, 571162624, 1438384149, 1587566, -668139240, 3, 921966},{131072, 0, 0, 1077575680, -1457127004, -443847898, 1256440772, 245366804, 1964032, -1787244896, 1073741825, 909791},{0, 0, 0, 807665664, -793074940, 627800, 226541568, 14, 1091267584, 1400882525, 403536600, 909613},{196608, 0, 0, 36077568, 408223923, 965779, -1223404472, 14, 2136469504, 222777925, 1470890006, 1120608},{0, 0, 0, 1175977984, -2143960454, 679272, -399310848, 55312402, 1344799, 2016739328, 1370488849, 1120543},{0, 35127296, 0, 1073741824, -1479212702, 1471328, 29332748, 17, -1819196416, -491029608, -725090293, 1531216},{0, 1, 0, 100663296, 1455587682, 1116820069, 1766479009, 2037645338, -1798391112, 632183157, -1695962987, 1386828},{0, 0, 0, -266076160, 1087750915, -1131850335, 1965609584, 18, -738197504, 567988877, 488112158, 611284},{131072, 16777264, 0, -469106688, -1252330125, -884192742, -500432215, 481675482, 1755926, 1580286336, 28, 1026048},{0, 16777216, 0, -1438941184, -788359051, 611288, 542446704, -1006108649, 1083346781, 1734612912, -1073741821, 1496127},{131072, 0, 0, -2046820352, -2143960659, 1220066, 257905824, 23, 1590272, 1409286144, -1019133224, 1523767},{0, 0, 0, 1141571584, -791534731, 1179602064, 686526040, -826691770, 1424716, -173064192, 22, 0},{262144, 83886080, 0, 402653184, -1587977468, 567378, -167772160, 19, -1043403776, 857327256, -714604517, 1595074},{196608, 0, 0, 33554432, 2041709197, -774720165, -280552127, -583008230, -725407832, -1916035948, -853278716, 1882324},{6144, 16777216, 0, 805306368, -192063476, -879923072, 727118465, -1894252532, -904752693, 130665668, -1933251185, 921876},{0, 0, 4096, 70942720, -425373813, 1037221264, -1359295295, -1814298621, 835785, -929803504, 1465705487, 254613},{0, 33554448, 0, -1607204576, -609620459, -1944953310, -196683543, -1955810342, -875487505, -1829729080, -859308014, 1767822},{0, 0, 0, 1378157920, -340614397, 428903844, 1397834184, -2147483639, 405808, -603979776, 1406926867, 1961430},{65536, 0, 0, 1513687648, 1957293572, 1762961965, 1255460137, -850564861, 232923, 0, 1570596544, 985607},{262144, 0, 4096, 1073741824, 31121986, -1677030613, 655378920, -2101084159, 1080435, -1275068416, 1240203292, 765702},{196608, 0, 8192, -2147483648, -1144970870, -732777114, -746238640, 11, 252117, -513206684, -702453482, 1136174},{0, 0, 0, 809041920, -1856626429, 1489568, -1729686552, 1, 773056512, -1075888123, 28, 248036},{0, 65, 0, -2143649792, -423550622, 1162646, 288266176, -1192391532, 1353233, 217864428, 1334837272, 921852},{0, 64, 0, 1881440256, 1102430469, -1752138351, -243526543, 906798935, 1582972650, 1956959753, -1719822582, 1132896},{0, 65, 0, -2146172928, 961717093, 611165, 1293883764, -243726461, 1557819263, 2030327648, -1722452400, 213399},{0, 0, -1342177280, 1111034112, -144872795, 814290, 1151827968, -917137519, 1119565, 228032512, -898629611, 1662119},{131072, 0, 0, 37290656, -640071262, 948952, -2025586688, -718975532, 1762729, 1342177280, 25, 1352704},{0, 64, 21256, 1077477376, -1529740956, -1777515286, -1788311192, -764057258, 1405736, 1811939328, -67120695, 1544723},{0, 48, 0, 805306368, 281698331, -1899452255, 1627050109, 46501137, 1669065, 0, 1492123648, 1081607},{0, 17, 0, -2046820352, 1510045836, 1489703, 134217728, 2008044868, 1975081, 1130239636, 378890077, 1516608},{0, 32, 0, 1882783744, 894607620, 1460783, -1216053248, 1492225628, -1325197435, 1095391472, 1221066775, 1440945},{0, 16777216, 0, 1744830464, 832676354, 678821, -196702608, -909563562, 264862, -681702932, 22, 1217536},{0, 18350080, 16384, 1646690304, 959512605, 1004125, 150769596, 264808335, -1483629374, 2139450412, -714037821, 1719913},{6144, 67108880, 0, -1321992192, -788088827, -1630628760, -1152584184, -1982736242, 5961568, 324984208, 14, 862367},{0, 64, 4096, 1547307328, -1178525684, 1226078, -1863499776, -2147483630, 1543921, -1527660544, -1893666420, 798504},{262336, 17825792, 0, 805306368, -614577902, -1064076382, 1876179599, -603081141, 826886345, -1160451755, 28, 1035264},{65536, 33554480, 0, -1073741824, -1710647214, -476992698, -1158686523, -1640746084, 1217264, -969719732, 12, 1926144},{2048, 0, 12288, 2359296, 117831680, -1026057081, -1019347475, -1037295860, 1807776, 765526576, -990380004, 612313},{0, 68206592, 128, -1342177280, -376524531, 705840602, -1945674307, 3, -623729664, 1590472459, -160356841, 1768334},{0, 0, 16520, 1174405120, -1496682830, 2144110050, -1197716000, -1073741796, -1085413951, -540405631, -1580219949, 1732433},{2048, 0, 16384, -1342177280, 1364845322, 798448681, 1332290520, 1073741837, 597049, 941244416, 1231590998, 773998},{0, 32, 0, 1880555520, 2018616069, 1338735725, -185984448, 1073741853, -288290064, 1770409732, 440500760, 650815},{0, 16777216, 16384, 100663296, 89842251, -1005490665, 1387530445, 1270449421, -2087187276, -1833297839, 1140898710, 1341380},{0, 16777216, 0, 1144684544, 2067098786, -863077291, -365625316, 1073741843, 1116213, -892564288, 1359508483, 1668479},{0, 16, 8192, -1841823744, -648621638, 1779334358, 1633145416, 116129815, 1859710808, -966781924, 356336207, 1316405},{0, 16777216, 8192, 808747008, 1755934738, 1481471467, 1275778025, -1051639999, 1472886608, 187585925, 1363673110, 1670823},{-2147483648, 64, 8192, 1077182464, -1464153181, -728777558, 632180048, -1345585131, -715884793, -1539092540, -2078738092, 1669699},{262144, 80, 4096, 1882753344, -70077942, 1758883036, 332668193, -1200881650, 1133463, 291542504, -663910826, 687766},{272576, 0, 1610612736, 2754208, 2008369408, -28418899, 1592015230, 1073741847, -1172777794, 1707842712, 17, 779264},{71680, 69730304, 0, -268140544, -1185496563, -1479707884, -1758924672, 1548222486, -1525647193, 1924411464, -668729333, 263621},{0, 0, 128, 805306368, 1899348748, 1124629593, 293913656, 11, 1523712, 4440064, 687079446, 1082255},{71680, 32, 0, 805306368, -70694630, -1747946078, -1304386447, -759845225, 1517380, -1757069300, -646343274, 1767659},{-2147483648, 17, 16384, 1879048192, -1051639779, 1489760, -1463546824, 1814366226, 1635205, -1456862140, 276299794, 183048},{0, 67633152, 0, -2076934144, -332826811, 2027000678, 1288887301, -1073741811, -1085673512, 1534049289, -684982248, 258424},{-2147479552, 50331712, 0, -1342177280, -631845348, -1324788520, -887493440, -1361262129, 934567, 787613940, -884998132, 990504},{65536, 64, 8192, 1174405120, -1413152603, 1473426, 167772160, -917766122, 922416, 222153540, 1265668060, 652215},{272448, 100663296, 0, 1882619904, 542794250, -266898799, 253014674, -633339882, 1633676, 2011404908, -1073741804, 1940562},{0, 67633152, 20480, -1342177280, -1875500532, 940696, 765509632, 1073741826, 1375859869, 2123726252, 167026449, 1177567},{0, 17, 16384, -268435456, -2143149291, 1199002, -923009024, -1610612721, -54314256, 2104039016, 312813120, 612921},{0, 0, 0, -1040187392, -506330453, 743148178, 794859352, -591563300, 650396, 492765888, -1030225892, 1446258},{0, 0, 8192, -2046820352, -1062641557, 1354706, 137576808, 3, -1845282816, -446428828, -1073741802, 1950269},{0, 67108880, 0, 1177092480, -1715906684, 1403436, 542284844, 1514259160, 911238, -901489768, 2, 1964032},{0, 0, 0, -1040187392, 1093772147, 1422355, -1768976108, 3, 1049982425, 1153143160, 1430116555, 1146199},{0, 0, 16384, 1107296256, -775519595, 1275280, 1171505152, -1933049827, 984983, 141843784, 1076205073, 1354293},{0, 64, 12288, 1142325248, -121976731, 566842390, -1001995176, 874268061, 1218437, -872415232, 356637842, 1853272},{0, 69730304, 0, -972488704, -786087542, 1058319256, 202408073, 1406664705, 686424, 257368064, 1247887183, 86027},{0, 0, 12288, -2113929216, 1439269450, -2112635479, 1143068761, 1469340738, 454211, 1568210944, -850068264, 1533505},{0, 0, 0, -2045214368, 1780556418, 1545771, 1145159680, 200918108, -1181348669, -1786323983, -1678720170, 1472980},{262144, 0, 0, 1142227296, 1549462666, 892073, -823079212, 417975247, 1140111, -453967872, -1673248693, 1045956},{0, 0, -2147483648, 103056800, -146388126, 1779674388, 223777200, -1789846782, 444726614, 1554501761, -952885028, 265498},{0, 0, 0, -2044100224, 1723924876, 780819051, 1099253369, -1073741801, 550206, 2092454892, -970671994, 1442883},{0, 0, 1746673664, 674508865, 2067614044, 1152359, -267691348, -626163071, 142404, 2082686028, -1072319719, 1859502},{0, 0, 16640, 37388576, -1506407518, 965740, -932456804, -1785652079, 1678519594, -2122934627, 1816492048, 1083057},{0, 0, 0, -2110420608, 1489663562, 642818909, -1943022355, -722730979, 423898159, 1447319436, -2077212268, 873920},{0, 0, -2011676672, 3672385, -80327936, 1289500, -1515191972, -674910203, 671926451, -1001011376, 1168397527, 960297},{262144, 0, 1207959552, 1144260032, 2067884707, 1146213, 238637100, 1265440792, 611646, 272203776, -1943528820, 1146993},{0, 67633152, -2013265920, -399209984, -356591534, 1175219366, 160373352, 68224463, 1151219721, -151913044, 119013399, 280646},{0, 67108880, -1879048192, 1714948640, -1230399422, 1461802, -241203928, -2147483639, -287567969, 1377799956, 1110503747, 1708114},{262144, 83886080, -1342177280, -2110125408, 734877827, -402093101, 236311140, 21, -1072674816, 1245254308, -830180975, 1480956},{393216, 16777216, 17024, 1141506048, 1788945235, 1808497571, -1499521620, -777995884, -1920809632, -234860128, -1218585827, 1387438},{0, 67108864, 0, -2076966624, -1137270411, 1538720, 1677721600, 9, 1612127232, 1849546524, -2093476087, 203922},{0, 0, 1344405504, 3836417, -709168640, 1277484, 603979776, 2, 1583135, 1438221400, 1146626652, 1599941},{0, 32, 0, -1073741824, -2133777582, -2058453990, -1917905600, 1366929181, 1500740, -729104384, 1219493911, 213373},{6144, 16, 0, 67108864, 388904004, -1018598635, 799285284, 58472028, 14547579, 1436012132, 1278787843, 1919206},{-2147483648, 67108865, 0, 1109983232, 1714875044, 1262931, 1094829168, 1610612757, 1406644, -1084751872, -638037426, 1233311},{0, 16, 0, -2076802816, -1253182875, 625582, -1275068416, -1073741824, -2087646704, 1353177185, 273707393, 1308038},{0, 0, 4096, -1342177280, 1104478733, 678491, 1514357788, 4, 1583362, 671088640, -954728432, 1952645},{0, 64, 0, 37126400, -1137540467, 621460, 805306368, 12, 992001, 0, -954662964, 1480961},{0, 0, 4096, 67108864, -1403600052, 1124881954, 1694472432, -1073741807, 1545965, -201326592, 119013391, 150257},{0, 16777216, 0, 70516736, -1404741469, -20359658, 1178960416, 28, 1157120, -232734208, -954728421, 475205},{0, 0, 0, -264568832, 1361453317, 808489, -2078146560, 11, 567395, 472154112, 1182540950, 1854324},{2048, 0, 0, 67108864, -1405762686, 1421934, 1796943776, 21, 0, -654671872, -2147483633, 1040497},{262144, 80, 0, 1107296256, -1043201452, 764754, -1082683496, -277348324, 1843006, 1090076672, 22, 464896},{131072, 16, 12288, 1879048192, -1674233758, -163033556, -1371356132, 26, 282112, 922140672, 1192755202, 1767159},{2048, 0, 0, 67108864, -1942677333, -195672540, -882252468, 17, 163840, -1527398400, -2147483643, 94321},{2048, 50331712, 0, -2080374784, -1405790035, 611886, -11608064, -1073741822, -208946494, -1827141820, 119013405, 1061108},{264192, 0, 0, 67108864, -1674394750, -326283730, -877645732, 12, -589838848, 1156337104, -1073741817, 465026},{0, 16777216, 0, -2144829440, -1405762749, 1005074, 1553252700, 9, -1824333824, -1682814640, 157324163, 1769569},{264384, 80, 0, 67108864, -1942147405, 76367406, -2042216901, 445644821, -1458309575, 1249139385, -2068840444, 94635},{65536, 67143248, 0, -1342177280, -1252659579, -993506456, -89143047, -672637607, 590335708, 1458666002, 460620557, 721349},{-1946157056, 100663362, 0, 1107296256, -1455095109, 611230, 1075167232, -223990654, 664619910, 304057384, 1277739286, 951844},{0, 81, 16512, -268435456, 1683835274, 1220139, 1209384960, 579872902, 780058, -1632630020, 687164683, 1885147},{201734208, 83886144, 8192, 1879048192, -1219577731, 655649364, 2131239903, -482677302, 266097, 1595670656, -775941988, 617257},{131072, 83904000, 16384, 1879048192, 1279965341, 938839, 638960228, 2, -2036334592, 1069900891, 1117529860, 1595946},{-2147155968, 16777281, 8192, 0, 917362688, 638485, 2142183772, 1039148505, 1782745, -695058432, 1104975639, 569886},{201601024, 83886193, 4096, 1879048192, 1546565717, -1110856147, 791322972, -480893620, 1951433271, 1189507152, -1644673972, 801421},{-2147155968, 100663360, 256, 1882783744, 1814485083, 588494357, -1895687524, 807936791, 541939544, 175391888, 1610612764, 1703746},{196608, 67108896, 21248, -1040187392, -1135683469, 1527316, 251724764, -1020240575, -4107715, -1752815804, 940048402, 839348},{262144, 50331648, 21256, 1073741824, -69885549, 1472038, 1443872768, 1083179017, 1351614719, 1584683648, 607852184, 1305271},{0, 87031808, 16768, -2113929216, 727040635, 695843, -1403174912, -1039565183, 449846816, -140056764, 1878006424, 986819},{0, 35127296, 16384, 1073741824, 741212555, 949803, -1409286144, -2147483637, 2051396793, 331659077, 148373519, 653154},{0, 83886144, 384, -2113929216, -1169800621, 1289758, 0, -1884815360, 1481469, -831238176, -274464753, 286490},{327680, 67158112, 28928, 1107296256, -1404741518, 1017384, -956850752, 1073741826, 1951883001, -165370242, -1348713399, 1446584},{0, 0, 0, 1073741824, -785800845, 1140964, 0, -1073741824, 1010945, 1157058588, 7, 1009664},{0, 0, 12288, -1073741824, -246029997, 1465890, 201326592, 8, 1006592, 1156157012, -2147483641, 1540852},{0, 0, 16768, 0, -1054768789, 943200, 0, 0, 1276065792, 1081365017, 889454607, 1146435},{137216, 83886144, 0, 0, 1277526403, -2096257507, -1507312244, 1073741829, 1670892, 1249132544, 1315700765, 969796},{0, 50331680, 0, 1073741824, -332291709, 685598, -534642688, 1073741826, 1147460, 841203712, 154787728, 94357},{0, 84934720, 12288, 1073741824, 2082578827, 1461781, -1872936960, 1149501443, -1484095976, -153274459, 1377304595, 1074000},{0, 0, 4096, -2080374784, 1548813130, 757275, -863825528, 13, 0, 644438656, 1158152219, 615340},{0, 67108880, 12288, 1140850688, 1547589796, 611869, -923598848, -1749286910, 1612354087, -1683249340, 255066134, 1068567},{0, 0, 16520, 1174405120, -1403406171, 611868, -299335024, 1073741847, 412967, -780337152, 1012012820, 1636016},{0, 16777216, 0, 1140850688, -62577758, 1405604, -1476395008, 26, -2087553707, 705729181, 1548484620, 149000},{0, 0, 0, 33554432, -1311153564, 888362, 0, 0, 708837376, 36291184, -2147483637, 94246},{0, 16777216, 0, 0, 473244276, 687657, 1543503872, 2, 499122176, -1030290972, 17, 600087},{0, 0, 0, 0, -2128281222, 868572, 1438777344, 2, 1795072, -1140850688, 81021713, 94401},{0, 0, 0, 1073741824, -1858264670, 868572, 0, -1073741824, 133196, -1946157056, 1519931972, 1744969},{0, 16777264, 0, 67108864, -1135208286, 806420, -872415232, 1163132951, 1069657, -78996628, 302629469, 779046},{71680, 0, 16640, 805306368, -870244340, -1496687070, 855814169, 131365634, 263231, 1749041152, 1693974545, 799490},{65536, 48, 8192, -1342177280, -1406281588, 1339313690, -568686596, -1073741821, 1048090, 188710912, 1517366424, 1054436},{196608, 0, 128, -2080374784, 407533669, 1087854107, -144502200, -2081423345, 1525069, 0, 605028352, 1738256},{131072, 50331648, 0, 1107296256, 2083879053, 636437, 238927872, 2, 0, -234881024, 54525967, 1569342},{0, 0, 4352, 0, 625124096, 1160751, -1509949440, 23, 0, 0, -536870912, 767673},{2048, 33554480, 0, 0, 0, 1397312, -621109248, 15, 1040896, -1509949440, 15, 0},{65536, 50331648, 256, 0, 0, 0, -1778384896, 15, 0, -1644167168, -536870897, 1951479},{-2147418112, 33554433, 0, 0, 0, 0, 1845493760, 1610612751, 1056503, 1778384896, 15, 0},{71680, 33554432, 0, 0, 0, 0, 1458954240, 14, 957952, 1241513984, 15, 0},{268288, 1, 4096, 0, 0, 0, -218914816, 536870941, 1379060, 0, 0, 1361408},{196608, 17825792, 0, 0, 0, 0, -973078528, 14, 0, 1861017992, 1073741838, 1937977},{0, 1572880, 8192, 0, 0, 0, 0, 0, 146944, -23781376, 29, 189952},{0, 32, 4096, 0, 0, 618688, 0, 0, 1735168, 167772160, 21, 1550848},{65536, 0, 8576, 0, 0, 0, -2113929216, 26, 0, -905969664, 536870938, 1150685},{69632, 0, 384, 0, 0, 0, -1104699392, 23, 0, 0, -536870912, 996908},{-2147483648, 1, 4352, 0, 0, 0, 0, 536870912, 1561421, 0, 1610612736, 167465},{0, 48, 4352, 0, 0, 0, 0, 0, 1220096, 1308622848, -536870884, 1748496},{-1946157056, 33554432, 0, 0, 0, 0, 0, 581304320, 171559, 1778384896, 2, 0},{-2013265920, 0, 12288, 0, 0, 0, 0, 1641938944, 619038, 0, 0, 156160},{0, 17825792, 12288, 0, 0, 0, 0, 0, 1162752, -675127296, 4, 154112},{2048, 33554432, 12288, 0, 0, 0, -1706237952, 26, 1140736, -1560150016, 26, 144896},{71680, 32, 0, 0, 0, 0, -1436983296, 20, 1844736, 0, 0, 1561088},{-2147352576, 0, 0, 0, 0, 1075392, -680247296, 1610612743, 1733184, 939524096, 22, 0},{6144, 16777248, 0, 0, 0, 0, 1176166400, 14, 1309184, 1912602624, 26, 0},{0, 0, 4096, 0, 0, 1400960, -637534208, 20, 0, 0, 0, 266752},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 254464},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, -1778384896, 3, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 1744830464, 17, 0, 0, 0, 1058816},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1327104, 0, 0, 0, 1073741824, 22, 1525760},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 548864, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1059840, 0, 0, 1141760},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 557056, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 1241513984, 23, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 1828929536, 17, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 813056, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 1275068416, 16, 1141760, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1089536, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 1811939328, 17, 1070080, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1343488, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 1543503872, 16, 1142784},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 548864, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 1879048192, 17, 1074176},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 802816, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1142784, -1946157056, 16, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1073152, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 1879048192, 17, 0, -1677721600, 16, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1335296, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, -1342177280, 16, 1143808},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 548864, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1098752, 1946157056, 17, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 819200, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1143808, -671088640, 16, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1073152, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 1946157056, 17, 0, -402653184, 16, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 1335296, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 1144832},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 565248, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1119232, 2013265920, 17, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 819200, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 1144832, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 524288, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{262144, 0, 0, 0, 0, 0, 2046820352, 17, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},{1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}};


//For 1st BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_A_addr;
reg [31:0]bram_ZYNQ_block_A_din;
wire [31:0]bram_ZYNQ_block_A_dout;
wire bram_ZYNQ_block_A_en;
wire [3:0]bram_ZYNQ_block_A_we;

//For 2nd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_B_addr;
reg [31:0]bram_ZYNQ_block_B_din;
wire [31:0]bram_ZYNQ_block_B_dout;
wire bram_ZYNQ_block_B_en;
wire [3:0]bram_ZYNQ_block_B_we;

//For 3rd BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_C_addr;
reg [31:0]bram_ZYNQ_block_C_din;
wire [31:0]bram_ZYNQ_block_C_dout;
wire bram_ZYNQ_block_C_en;
wire [3:0]bram_ZYNQ_block_C_we;

//For 4th BRAM
wire [ADDR_WIDTH_DATA_BRAM - 1 : 0]bram_ZYNQ_block_D_addr;
reg [31:0]bram_ZYNQ_block_D_din;
wire [31:0]bram_ZYNQ_block_D_dout;
wire bram_ZYNQ_block_D_en;
wire [3:0]bram_ZYNQ_block_D_we;

//Instruction BRAM
wire [31:0]bram_ZYNQ_INST_addr;
wire bram_ZYNQ_INST_en;
wire bram_ZYNQ_INST_we;

wire [31:0]bram_ZYNQ_INST_din_part_0;
wire [31:0]bram_ZYNQ_INST_din_part_1;
wire [31:0]bram_ZYNQ_INST_din_part_2;
wire [31:0]bram_ZYNQ_INST_din_part_3;
wire [31:0]bram_ZYNQ_INST_din_part_4;
wire [31:0]bram_ZYNQ_INST_din_part_5;
wire [31:0]bram_ZYNQ_INST_din_part_6;
wire [31:0]bram_ZYNQ_INST_din_part_7;
wire [31:0]bram_ZYNQ_INST_din_part_8;
wire [31:0]bram_ZYNQ_INST_din_part_9;
wire [31:0]bram_ZYNQ_INST_din_part_10;
wire [31:0]bram_ZYNQ_INST_din_part_11;

wire [31:0]bram_ZYNQ_INST_dout_part_0;
wire [31:0]bram_ZYNQ_INST_dout_part_1;
wire [31:0]bram_ZYNQ_INST_dout_part_2;
wire [31:0]bram_ZYNQ_INST_dout_part_3;
wire [31:0]bram_ZYNQ_INST_dout_part_4;
wire [31:0]bram_ZYNQ_INST_dout_part_5;
wire [31:0]bram_ZYNQ_INST_dout_part_6;
wire [31:0]bram_ZYNQ_INST_dout_part_7;
wire [31:0]bram_ZYNQ_INST_dout_part_8;
wire [31:0]bram_ZYNQ_INST_dout_part_9;
wire [31:0]bram_ZYNQ_INST_dout_part_10;
wire [31:0]bram_ZYNQ_INST_dout_part_11;

//debug signals
wire [1:0]debug_state;

reg [31:0]BRAM_dump[0:3][0:2047];
reg [31:0]fptr,fptr2;
integer count;
reg complete_bit;

//Mux signals
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_A_dout;
reg [1:0]sel_mux_dataBRAM;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_B_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_C_dout;

reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_0; //For dumping BRAM contents
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_1; //For clearing
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_2; //For loading A matrix
reg [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_3; //Currently unused
wire [ADDR_WIDTH_DATA_BRAM-1:0]mux_dataBRAM_D_dout;

reg mux_dataBRAM_A_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_en1 = 0; //For clearing
reg mux_dataBRAM_A_en2 = 0; //For loading A matrix
reg mux_dataBRAM_A_en3 = 0; //Currently unused
wire mux_dataBRAM_A_endout;

reg mux_dataBRAM_B_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_en1 = 0; //For clearing
reg mux_dataBRAM_B_en2 = 0; //For loading A matrix
reg mux_dataBRAM_B_en3 = 0; //Currently unused
wire mux_dataBRAM_B_endout;

reg mux_dataBRAM_C_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_en1 = 0; //For clearing
reg mux_dataBRAM_C_en2 = 0; //For loading A matrix
reg mux_dataBRAM_C_en3 = 0; //Currently unused
wire mux_dataBRAM_C_endout;

reg mux_dataBRAM_D_en0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_en1 = 0; //For clearing
reg mux_dataBRAM_D_en2 = 0; //For loading A matrix
reg mux_dataBRAM_D_en3 = 0; //Currently unused
wire mux_dataBRAM_D_endout;

reg mux_dataBRAM_A_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_A_we1 = 0; //For clearing
reg mux_dataBRAM_A_we2 = 0; //For loading A matrix
reg mux_dataBRAM_A_we3 = 0; //Currently unused
wire mux_dataBRAM_A_wedout;

reg mux_dataBRAM_B_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_B_we1 = 0; //For clearing
reg mux_dataBRAM_B_we2 = 0; //For loading A matrix
reg mux_dataBRAM_B_we3 = 0; //Currently unused
wire mux_dataBRAM_B_wedout;

reg mux_dataBRAM_C_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_C_we1 = 0; //For clearing
reg mux_dataBRAM_C_we2 = 0; //For loading A matrix
reg mux_dataBRAM_C_we3 = 0; //Currently unused
wire mux_dataBRAM_C_wedout;

reg mux_dataBRAM_D_we0 = 0; //For dumping BRAM contents
reg mux_dataBRAM_D_we1 = 0; //For clearing
reg mux_dataBRAM_D_we2 = 0; //For loading A matrix
reg mux_dataBRAM_D_we3 = 0; //Currently unused
wire mux_dataBRAM_D_wedout;

reg [31:0]mux_dataBRAM_A_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_A_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_A_din_out;
reg sel_mux_dataBRAM_din;

reg [31:0]mux_dataBRAM_B_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_B_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_B_din_out;

reg [31:0]mux_dataBRAM_C_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_C_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_C_din_out;

reg [31:0]mux_dataBRAM_D_din0; //for clearing the data BRAMS
reg [31:0]mux_dataBRAM_D_din1; //for loading the data BRAMS
wire [31:0]mux_dataBRAM_D_din_out;

//Instruction BRAM muxes
reg [31:0]instBRAM_part0_din;
reg [31:0]instBRAM_part1_din;
reg [31:0]instBRAM_part2_din;
reg [31:0]instBRAM_part3_din;
reg [31:0]instBRAM_part4_din;
reg [31:0]instBRAM_part5_din;
reg [31:0]instBRAM_part6_din;
reg [31:0]instBRAM_part7_din;
reg [31:0]instBRAM_part8_din;
reg [31:0]instBRAM_part9_din;
reg [31:0]instBRAM_part10_din;
reg [31:0]instBRAM_part11_din;

reg instBRAM_en = 0;
reg instBRAM_we = 0;
reg [ADDR_WIDTH-1:0]instBRAM_addr;


//Memory dump start and complete signals
reg start_mem_dump;
reg mem_dump_complete;
reg start_dataBRAM_erase;
reg dataBRAM_erase_complete;
reg start_A_load;
reg A_load_complete;
reg start_instBRAM_erase;
reg instBRAM_erase_complete;
reg start_inst_load;
reg inst_load_complete;
reg start_full_run;
reg complete_full_run;
reg start0; //For full run
reg complete_sig;

LUDH_TEST_WRAPPER #(ADDR_WIDTH,ADDR_WIDTH_DATA_BRAM,CTRL_WIDTH,AU_SEL_WIDTH,BRAM_SEL_WIDTH) uut1 (
CLK_100,
CLK_200,
locked,
RST_IN,
start_sig,
completed,

//First BRAM
bram_ZYNQ_block_A_addr, 
bram_ZYNQ_block_A_din, 
bram_ZYNQ_block_A_dout, 
bram_ZYNQ_block_A_en,
bram_ZYNQ_block_A_we, 

//Second BRAM
bram_ZYNQ_block_B_addr, 
bram_ZYNQ_block_B_din, 
bram_ZYNQ_block_B_dout, 
bram_ZYNQ_block_B_en,
bram_ZYNQ_block_B_we, 

//Third BRAM
bram_ZYNQ_block_C_addr, 
bram_ZYNQ_block_C_din, 
bram_ZYNQ_block_C_dout, 
bram_ZYNQ_block_C_en,
bram_ZYNQ_block_C_we, 

//Fourth BRAM
bram_ZYNQ_block_D_addr, 
bram_ZYNQ_block_D_din, 
bram_ZYNQ_block_D_dout, 
bram_ZYNQ_block_D_en,
bram_ZYNQ_block_D_we, 

//Instruction BRAM
bram_ZYNQ_INST_addr,
bram_ZYNQ_INST_en,
bram_ZYNQ_INST_we,
        
bram_ZYNQ_INST_din_part_0,
bram_ZYNQ_INST_din_part_1,
bram_ZYNQ_INST_din_part_2,
bram_ZYNQ_INST_din_part_3,
bram_ZYNQ_INST_din_part_4,
bram_ZYNQ_INST_din_part_5,
bram_ZYNQ_INST_din_part_6,
bram_ZYNQ_INST_din_part_7,
bram_ZYNQ_INST_din_part_8,
bram_ZYNQ_INST_din_part_9,
bram_ZYNQ_INST_din_part_10,
bram_ZYNQ_INST_din_part_11,
        
bram_ZYNQ_INST_dout_part_0,
bram_ZYNQ_INST_dout_part_1,
bram_ZYNQ_INST_dout_part_2,
bram_ZYNQ_INST_dout_part_3,
bram_ZYNQ_INST_dout_part_4,
bram_ZYNQ_INST_dout_part_5,
bram_ZYNQ_INST_dout_part_6,
bram_ZYNQ_INST_dout_part_7,
bram_ZYNQ_INST_dout_part_8,
bram_ZYNQ_INST_dout_part_9,
bram_ZYNQ_INST_dout_part_10,
bram_ZYNQ_INST_dout_part_11,
        
//debug signals
debug_state
);

initial begin
CLK_100 = 1'b1;
forever #(t_100/2) CLK_100 = ~CLK_100;
end

initial begin
CLK_200 = 1'b1;
forever #(t_200/2) CLK_200 = ~CLK_200;
end

//Initiallizing the mux to be used for DATA BRAMS address multiplexing
//For address
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut2(mux_dataBRAM_A_dout,mux_dataBRAM_A_0,mux_dataBRAM_A_1,mux_dataBRAM_A_2,mux_dataBRAM_A_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut3(mux_dataBRAM_B_dout,mux_dataBRAM_B_0,mux_dataBRAM_B_1,mux_dataBRAM_B_2,mux_dataBRAM_B_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut4(mux_dataBRAM_C_dout,mux_dataBRAM_C_0,mux_dataBRAM_C_1,mux_dataBRAM_C_2,mux_dataBRAM_C_3,sel_mux_dataBRAM);
mux_4x1 #(ADDR_WIDTH_DATA_BRAM) uut5(mux_dataBRAM_D_dout,mux_dataBRAM_D_0,mux_dataBRAM_D_1,mux_dataBRAM_D_2,mux_dataBRAM_D_3,sel_mux_dataBRAM);

//For enable
mux_4x1 #(1) uut6(mux_dataBRAM_A_endout,mux_dataBRAM_A_en0,mux_dataBRAM_A_en1,mux_dataBRAM_A_en2,mux_dataBRAM_A_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut7(mux_dataBRAM_B_endout,mux_dataBRAM_B_en0,mux_dataBRAM_B_en1,mux_dataBRAM_B_en2,mux_dataBRAM_B_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut8(mux_dataBRAM_C_endout,mux_dataBRAM_C_en0,mux_dataBRAM_C_en1,mux_dataBRAM_C_en2,mux_dataBRAM_C_en3,sel_mux_dataBRAM);
mux_4x1 #(1) uut9(mux_dataBRAM_D_endout,mux_dataBRAM_D_en0,mux_dataBRAM_D_en1,mux_dataBRAM_D_en2,mux_dataBRAM_D_en3,sel_mux_dataBRAM);

//For Write enable
mux_4x1 #(1) uut10(mux_dataBRAM_A_wedout,mux_dataBRAM_A_we0,mux_dataBRAM_A_we1,mux_dataBRAM_A_we2,mux_dataBRAM_A_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut11(mux_dataBRAM_B_wedout,mux_dataBRAM_B_we0,mux_dataBRAM_B_we1,mux_dataBRAM_B_we2,mux_dataBRAM_B_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut12(mux_dataBRAM_C_wedout,mux_dataBRAM_C_we0,mux_dataBRAM_C_we1,mux_dataBRAM_C_we2,mux_dataBRAM_C_we3,sel_mux_dataBRAM);
mux_4x1 #(1) uut13(mux_dataBRAM_D_wedout,mux_dataBRAM_D_we0,mux_dataBRAM_D_we1,mux_dataBRAM_D_we2,mux_dataBRAM_D_we3,sel_mux_dataBRAM);

//For din
mux_2x1 #(32) uut14(mux_dataBRAM_A_din_out,mux_dataBRAM_A_din0,mux_dataBRAM_A_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut15(mux_dataBRAM_B_din_out,mux_dataBRAM_B_din0,mux_dataBRAM_B_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut16(mux_dataBRAM_C_din_out,mux_dataBRAM_C_din0,mux_dataBRAM_C_din1,sel_mux_dataBRAM_din);
mux_2x1 #(32) uut17(mux_dataBRAM_D_din_out,mux_dataBRAM_D_din0,mux_dataBRAM_D_din1,sel_mux_dataBRAM_din);


initial begin
start_mem_dump <= 0;
mem_dump_complete <= 0;
start_dataBRAM_erase <= 0;
dataBRAM_erase_complete <= 0;
start_A_load <= 0;
A_load_complete <= 0;
start_instBRAM_erase <= 0;
instBRAM_erase_complete <= 0;
start_inst_load <= 0;
inst_load_complete <= 0;
complete_full_run <= 0;
sel_mux_dataBRAM <= 2'b00;
sel_mux_dataBRAM_din <= 1'b0;

count <= -1;
complete_bit <= 1'b0;
locked <= 1'b0;

#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
RST_IN <= 1'b1;

//Resetting the contents of data BRAMS and Inst BRAM
#(t_100*50)
sel_mux_dataBRAM <= 2'b01;
sel_mux_dataBRAM_din <= 1'b0;
start_dataBRAM_erase <= 1'b1;

@(posedge dataBRAM_erase_complete)
#(t_100*50)
start_dataBRAM_erase <= 0;

#(t_100*50)
start_instBRAM_erase <= 1'b1;

@(posedge instBRAM_erase_complete)
#(t_100*50)
start_instBRAM_erase <= 0;

//Loading the A matrix
#(t_100*50)
sel_mux_dataBRAM <= 2'b10;
sel_mux_dataBRAM_din <= 1'b1;
start_A_load <= 1'b1;

@(posedge A_load_complete)
#(t_100*50)
start_A_load <= 0;

//RST = 0
#(t_100*50)
RST_IN <= 1'b0;

//Locked = 1
#(t_100*50)
locked <= 1'b1;

//Loading the instruction matrix and starting LU Decomposition
#(t_100*50)
start_full_run = 1'b1;

@(posedge complete_sig)
complete_bit <= 1'b1;
#(t_100*50)
start_full_run <= 1'b0;

#(t_100*50)
sel_mux_dataBRAM <= 2'b00;
start_mem_dump <= 1;

@(posedge mem_dump_complete)
#(t_100*50)
start_mem_dump <= 0;
$stop;

end

assign start_sig = start0;
assign complete_sig = complete_full_run;

//Address signals(data BRAM)
assign bram_ZYNQ_block_A_addr = mux_dataBRAM_A_dout;
assign bram_ZYNQ_block_B_addr = mux_dataBRAM_B_dout;
assign bram_ZYNQ_block_C_addr = mux_dataBRAM_C_dout;
assign bram_ZYNQ_block_D_addr = mux_dataBRAM_D_dout;

//Enable signals(data BRAM)
assign bram_ZYNQ_block_A_en = mux_dataBRAM_A_endout;
assign bram_ZYNQ_block_B_en = mux_dataBRAM_B_endout;
assign bram_ZYNQ_block_C_en = mux_dataBRAM_C_endout;
assign bram_ZYNQ_block_D_en = mux_dataBRAM_D_endout;

//Write enable signals(data BRAM)
assign bram_ZYNQ_block_A_we = mux_dataBRAM_A_wedout;
assign bram_ZYNQ_block_B_we = mux_dataBRAM_B_wedout;
assign bram_ZYNQ_block_C_we = mux_dataBRAM_C_wedout;
assign bram_ZYNQ_block_D_we = mux_dataBRAM_D_wedout;

//din signals(data BRAM)
assign bram_ZYNQ_block_A_din = mux_dataBRAM_A_din_out;
assign bram_ZYNQ_block_B_din = mux_dataBRAM_B_din_out;
assign bram_ZYNQ_block_C_din = mux_dataBRAM_C_din_out;
assign bram_ZYNQ_block_D_din = mux_dataBRAM_D_din_out;

//Address signal(inst BRAM)
assign bram_ZYNQ_INST_addr = instBRAM_addr;

//Enable signal(inst BRAM)
assign bram_ZYNQ_INST_en = instBRAM_en;

//Write enable signal(inst BRAM)
assign bram_ZYNQ_INST_we = instBRAM_we;

//din signal(inst BRAM)
assign bram_ZYNQ_INST_din_part_0 = instBRAM_part0_din;
assign bram_ZYNQ_INST_din_part_1 = instBRAM_part1_din;
assign bram_ZYNQ_INST_din_part_2 = instBRAM_part2_din;
assign bram_ZYNQ_INST_din_part_3 = instBRAM_part3_din;
assign bram_ZYNQ_INST_din_part_4 = instBRAM_part4_din;
assign bram_ZYNQ_INST_din_part_5 = instBRAM_part5_din;
assign bram_ZYNQ_INST_din_part_6 = instBRAM_part6_din;
assign bram_ZYNQ_INST_din_part_7 = instBRAM_part7_din;
assign bram_ZYNQ_INST_din_part_8 = instBRAM_part8_din;
assign bram_ZYNQ_INST_din_part_9 = instBRAM_part9_din;
assign bram_ZYNQ_INST_din_part_10 = instBRAM_part10_din;
assign bram_ZYNQ_INST_din_part_11 = instBRAM_part11_din;


//Always block for full run
always@(posedge CLK_100) begin
if(CLK_100  == 1 && start_full_run == 1 && complete_full_run != 1) begin
//Start loading complete instructions
start_inst_load <= 1'b1;
@(posedge inst_load_complete)
#(t_100*50)
start_inst_load <= 0;

//Start the LU Decomposition
#(t_100*50)
start0 <= 1'b1;
complete_full_run <= 1'b0;

//Waiting for completion
@(posedge completed)
complete_full_run <= 1'b1;

end
else if(CLK_100 == 1 && start_full_run == 0) begin
start0 <= 0;
complete_full_run <= 0;
end
end

//Always block to dump bram contents
always@(posedge CLK_200) begin
if(CLK_200 == 1 && start_mem_dump == 1 && mem_dump_complete != 1)begin 

    if(count == -1) begin
        fptr = $fopen("BRAM_dump.txt","w");
        $fdisplay(fptr,"float bram_dump[%d][%d];",4,2**ADDR_WIDTH_DATA_BRAM);
        mux_dataBRAM_A_en0 = 1'b1; mux_dataBRAM_B_en0 = 1'b1; mux_dataBRAM_C_en0 = 1'b1; mux_dataBRAM_D_en0 = 1'b1;
        mux_dataBRAM_A_we0 = 1'b0; mux_dataBRAM_B_we0 = 1'b0; mux_dataBRAM_C_we0 = 1'b0; mux_dataBRAM_D_we0 = 1'b0;
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];
    end
    else if(count == 0) begin
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Addres
    end
    else if(count <= 2048 && count >= 1)begin
        $fdisplay(fptr,"bram_dump[0][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_A_dout)); //count-1 because BRAM has single cycle latency
        $fdisplay(fptr,"bram_dump[1][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_B_dout));
        $fdisplay(fptr,"bram_dump[2][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_C_dout));
        $fdisplay(fptr,"bram_dump[3][%d] = %e;",count-1,float_conv(bram_ZYNQ_block_D_dout));
        count = count + 1;
        mux_dataBRAM_A_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_0 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_0 = count[ADDR_WIDTH_DATA_BRAM-1:0];//Address
    end
    else if (count == 2049) begin
        $fclose(fptr);
        count = -1;
        mem_dump_complete = 1;    
        mux_dataBRAM_A_en0 = 1'b0; mux_dataBRAM_B_en0 = 1'b0; mux_dataBRAM_C_en0 = 1'b0; mux_dataBRAM_D_en0 = 1'b0;   
    end
end
else if(CLK_200 == 1 && start_mem_dump == 0)
    mem_dump_complete = 0;
end


//Always block to erase data BRAM contents
always@(posedge CLK_200) begin
if(CLK_200 == 1 && start_dataBRAM_erase == 1 && dataBRAM_erase_complete != 1)begin 

    if(count <= 2048-2 && count >= -1)begin
        if(count == -1) begin
            mux_dataBRAM_A_en1 = 1'b1; mux_dataBRAM_B_en1 = 1'b1; mux_dataBRAM_C_en1 = 1'b1; mux_dataBRAM_D_en1 = 1'b1;
            mux_dataBRAM_A_we1 = 1'b1; mux_dataBRAM_B_we1 = 1'b1; mux_dataBRAM_C_we1 = 1'b1; mux_dataBRAM_D_we1 = 1'b1;
            mux_dataBRAM_A_din0 = 0; mux_dataBRAM_B_din0 = 0; mux_dataBRAM_C_din0 = 0; mux_dataBRAM_D_din0 = 0; //Reset value
        end
        count = count + 1;
        mux_dataBRAM_A_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_B_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_C_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; mux_dataBRAM_D_1 = count[ADDR_WIDTH_DATA_BRAM-1:0]; //Address
    end
    else if (count == 2048-1) begin
        count = -1;
        dataBRAM_erase_complete = 1;   
        mux_dataBRAM_A_en1 = 1'b0; mux_dataBRAM_B_en1 = 1'b0; mux_dataBRAM_C_en1 = 1'b0; mux_dataBRAM_D_en1 = 1'b0;
        mux_dataBRAM_A_we1 = 1'b0; mux_dataBRAM_B_we1 = 1'b0; mux_dataBRAM_C_we1 = 1'b0; mux_dataBRAM_D_we1 = 1'b0;    
    end
end
else if(CLK_200 == 1 && start_dataBRAM_erase == 0)
    dataBRAM_erase_complete = 0;
end

//Always block to load the A matrix in data bram
always@(posedge CLK_200) begin
if(CLK_200 == 1 && start_A_load == 1 && A_load_complete != 1)begin 

    if(count <= A_size-2 && count >= -1)begin
        if(count == -1) //Initialization of en signals
            mux_dataBRAM_A_en2 = 1'b1; mux_dataBRAM_B_en2 = 1'b1; mux_dataBRAM_C_en2 = 1'b1; mux_dataBRAM_D_en2 = 1'b1;
            
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0;//Initially assigning all the write enables to 0
        count = count + 1;
        if(A_BRAMInd[count] == 0) begin//making one of the write enables 1
            mux_dataBRAM_A_we2 = 1'b1; mux_dataBRAM_A_2 = A_BRAMAddr[count]; mux_dataBRAM_A_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 1) begin
            mux_dataBRAM_B_we2 = 1'b1; mux_dataBRAM_B_2 = A_BRAMAddr[count]; mux_dataBRAM_B_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 2) begin
            mux_dataBRAM_C_we2 = 1'b1; mux_dataBRAM_C_2 = A_BRAMAddr[count]; mux_dataBRAM_C_din1 = A[count];
        end
        else if(A_BRAMInd[count] == 3) begin
            mux_dataBRAM_D_we2 = 1'b1; mux_dataBRAM_D_2 = A_BRAMAddr[count]; mux_dataBRAM_D_din1 = A[count];
        end
    end
    else if (count == A_size-1) begin
        count = -1;
        A_load_complete = 1;   
        mux_dataBRAM_A_en2 = 1'b0; mux_dataBRAM_B_en2 = 1'b0; mux_dataBRAM_C_en2 = 1'b0; mux_dataBRAM_D_en2 = 1'b0;
        mux_dataBRAM_A_we2 = 1'b0; mux_dataBRAM_B_we2 = 1'b0; mux_dataBRAM_C_we2 = 1'b0; mux_dataBRAM_D_we2 = 1'b0;    
    end
end
else if(CLK_200 == 1 && start_A_load == 0)
    A_load_complete = 0;
end

//Always block to erase inst BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_instBRAM_erase == 1 && instBRAM_erase_complete != 1)begin 

    if(count <= 4096-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
            instBRAM_part0_din = 0; instBRAM_part1_din = 0; instBRAM_part2_din = 0; instBRAM_part3_din = 0; instBRAM_part4_din = 0; instBRAM_part5_din = 0;
            instBRAM_part6_din = 0; instBRAM_part7_din = 0; instBRAM_part8_din = 0; instBRAM_part9_din = 0; instBRAM_part10_din = 0; instBRAM_part11_din = 0;
        end
        count = count + 1;
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == 4096-1) begin
        count = -1;
        instBRAM_erase_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_instBRAM_erase == 0)
    instBRAM_erase_complete = 0;
end

//Always block to load instruction to instruction BRAM
always@(posedge CLK_100) begin
if(CLK_100 == 1 && start_inst_load == 1 && inst_load_complete != 1)begin 

    if(count <= total_instructions-2 && count >= -1)begin
        if(count == -1) begin
            instBRAM_en = 1'b1;
            instBRAM_we = 1'b1;
        end
        count = count + 1;
        instBRAM_part0_din = Inst[count][0]; instBRAM_part1_din = Inst[count][1]; instBRAM_part2_din = Inst[count][2]; instBRAM_part3_din = Inst[count][3]; 
        instBRAM_part4_din = Inst[count][4]; instBRAM_part5_din = Inst[count][5]; instBRAM_part6_din = Inst[count][6]; instBRAM_part7_din = Inst[count][7]; 
        instBRAM_part8_din = Inst[count][8]; instBRAM_part9_din = Inst[count][9]; instBRAM_part10_din = Inst[count][10]; instBRAM_part11_din = Inst[count][11];
        instBRAM_addr = count[ADDR_WIDTH-1:0];
    end
    else if (count == total_instructions-1) begin
        count = -1;
        inst_load_complete = 1;   
        instBRAM_en = 1'b0;
        instBRAM_we = 1'b0;
    end
end
else if(CLK_100 == 1 && start_inst_load == 0)
    inst_load_complete = 0;
end

function real float_conv(input [31:0]b_num);
reg sign;
reg [7:0]weighted_expt;
integer actual_expt;
reg [1:23] mantissa;
reg [7:0] i;
real temp_result,temp_decimal;

begin
sign = b_num >> 31;
weighted_expt = (b_num & 32'h7f800000)>> 23;
mantissa = b_num & 32'h007fffff;

if(weighted_expt == 0)begin
	temp_result = 1.0;
	for(i=0;i<126;i=i+1)
		temp_result = temp_result/2;

	temp_decimal = 0;
	for(i=1;i<=23;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(1.0/(1<<i));
		
	temp_result = temp_result*temp_decimal;
	if(sign==1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
	end
else if(weighted_expt>0 && weighted_expt <255) begin
	actual_expt = weighted_expt-127;
	if(actual_expt<0)begin
		temp_result = 1.0;
		actual_expt = -actual_expt;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result/2;
		end
	else begin
		temp_result = 1.0;
		for(i=0;i<actual_expt;i=i+1)
			temp_result = temp_result*2;
	end

	temp_decimal = 0;
	for(i=1;i<=23;i=i+1)
		temp_decimal = temp_decimal + mantissa[i]*(1.0/(1<<i));

	temp_decimal = temp_decimal + 1;
	temp_result = temp_result*temp_decimal;
	if(sign == 1)
		float_conv = -temp_result;
	else
		float_conv = temp_result;
end
else if(weighted_expt == 255)begin
/*if(mantissa == 0 and sign == 0)
float_conv = "inf";
else if(mantissa == 0 and sign == 1)
float_conv = "-inf";
else
float_conv = "nan";*/
end

end
endfunction

endmodule

module mux_4x1 #(parameter integer data_width = 11)(dout,din0,din1,din2,din3,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input [data_width-1:0]din2;
input [data_width-1:0]din3;
input [1:0]sel;

always@(din0,din1,din2,din3,sel) begin
case(sel)
2'b00: dout <= din0;
2'b01: dout <= din1;
2'b10: dout <= din2;
2'b11: dout <= din3;
endcase
end
endmodule

module mux_2x1 #(parameter integer data_width = 32)(dout,din0,din1,sel);
output reg [data_width-1:0]dout;
input [data_width-1:0]din0;
input [data_width-1:0]din1;
input sel;

always@(din0,din1,sel) begin
case(sel)
1'b0: dout <= din0;
1'b1: dout <= din1;
endcase
end
endmodule













